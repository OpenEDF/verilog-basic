module hello_pli;
    
initial begin
   $hello;
   #20 $finish;
end

endmodule
