package router_stimulus_pkg;

import uvm_pkg::*;

`include "packet.sv"

// Lab 2: Task 8, Step 2 - include the packet_sequence.sv file
//
// ToDo
`include "packet_sequence.sv"



// Lab 2: Task 10, Step 2 - include the packet_da_3.sv file
//
// ToDo
`include "packet_da_3.sv"



endpackage
