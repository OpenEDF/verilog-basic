//
// Book, "RTL Modeling with SystemVerilog for ASIC and FPGA Design"
// by Stuart Sutherland
//
// N-bit 2:1 multiplexor modeled with an if-else statement.
//
// Copyright 2016, Stuart Sutherland. All rights reserved.
//
// Version 1.0
//

`begin_keywords "1800-2012" // use SystemVerilog-2012 keywords
module mux2to1
#(parameter N = 4)            // bus size
(input  logic         sel,    // 1-bit input
 input  logic [N-1:0] a, b,   // scalable input size
 output logic [N-1:0] y       // scalable output size
);
  timeunit 1ns/1ns;

  always_comb begin
    if (sel) y = a; 
    else     y = b;
  end

endmodule: mux2to1
`end_keywords
