/**********************************************************************
 * Using enumerated type methods to print label names
 *
 * Author: Stuart Sutherland
 *
 * (c) Copyright 2003, Sutherland HDL, Inc. *** ALL RIGHTS RESERVED ***
 * www.sutherland-hdl.com
 *
 * Used with permission in the book, "SystemVerilog for Design"
 *  By Stuart Sutherland, Simon Davidmann, and Peter Flake.
 *  Book copyright: 2003, Kluwer Academic Publishers, Norwell, MA, USA
 *  www.wkap.il, ISBN: 0-4020-7530-8
 *
 * Revision History:
 *   1.00 15 Dec 2003 -- original code, as included in book
 *   1.01 10 Jul 2004 -- cleaned up comments, added expected results
 *                       to output messages
 *
 * Caveat: Expected results displayed for this code example are based
 * on an interpretation of the SystemVerilog 3.1 standard by the code
 * author or authors.  At the time of writing, official SystemVerilog
 * validation suites were not available to validate the example.
 *
 * RIGHT TO USE: This code example, or any portion thereof, may be
 * used and distributed without restriction, provided that this entire
 * comment block is included with the example.
 *
 * DISCLAIMER: THIS CODE EXAMPLE IS PROVIDED "AS IS" WITHOUT WARRANTY
 * OF ANY KIND, EITHER EXPRESS OR IMPLIED, INCLUDING, BUT NOT LIMITED
 * TO WARRANTIES OF MERCHANTABILITY, FITNESS OR CORRECTNESS. IN NO
 * EVENT SHALL THE AUTHOR OR AUTHORS BE LIABLE FOR ANY DAMAGES,
 * INCLUDING INCIDENTAL OR CONSEQUENTIAL DAMAGES, ARISING OUT OF THE
 * USE OF THIS CODE.
 *********************************************************************/

module FSM (input wire resetN, clock);

  enum bit [1:0] {WAITE=2'b01, LOAD=2'b10, READY} State, Next;

  always @(posedge clock, negedge resetN)
    if (!resetN) State <= READY;
    else         State <= Next;

  always @(State)
    begin
      $display("\nCurrent state is %s (%b)", State.name, State);
      case (State)
        WAITE: Next = LOAD;
        LOAD:  Next = READY;
        READY: Next = WAITE;
      endcase
      $display("Next state will be %s (%b)", Next.name, Next);
    end
endmodule


module test;

  logic clock, resetN;

  FSM dut (.clock(clock), .resetN(resetN) );

  initial begin
    clock = 0;
    forever #5 clock = ~clock;
  end

  initial begin
    $display("\n Expect State to sequence through READY, WAITE, LOAD, READY");
    $display(" Expect Next to sequence through WAITE, LOAD, READY, WAITE\n");
    resetN <= 0;
    #8 resetN =1;
    repeat(4) @(negedge clock) ;
    $display("");
    $finish;
  end

endmodule
