/**********************************************************************
 * Restrictions on  passing unpacked structures through module ports
 * (must be declared with same typedef on both sides of port)
 *
 * Author: Stuart Sutherland
 *
 * (c) Copyright 2003, Sutherland HDL, Inc. *** ALL RIGHTS RESERVED ***
 * www.sutherland-hdl.com
 *
 * Used with permission in the book, "SystemVerilog for Design"
 *  By Stuart Sutherland, Simon Davidmann, and Peter Flake.
 *  Book copyright: 2003, Kluwer Academic Publishers, Norwell, MA, USA
 *  www.wkap.il, ISBN: 0-4020-7530-8
 *
 * Revision History:
 *   1.00 15 Dec 2003 -- original code, as included in book
 *   1.01 10 Jul 2004 -- cleaned up comments, added expected results
 *                       to output messages
 *
 * Caveat: Expected results displayed for this code example are based
 * on an interpretation of the SystemVerilog 3.1 standard by the code
 * author or authors.  At the time of writing, official SystemVerilog
 * validation suites were not available to validate the example.
 *
 * RIGHT TO USE: This code example, or any portion thereof, may be
 * used and distributed without restriction, provided that this entire
 * comment block is included with the example.
 *
 * DISCLAIMER: THIS CODE EXAMPLE IS PROVIDED "AS IS" WITHOUT WARRANTY
 * OF ANY KIND, EITHER EXPRESS OR IMPLIED, INCLUDING, BUT NOT LIMITED
 * TO WARRANTIES OF MERCHANTABILITY, FITNESS OR CORRECTNESS. IN NO
 * EVENT SHALL THE AUTHOR OR AUTHORS BE LIABLE FOR ANY DAMAGES,
 * INCLUDING INCIDENTAL OR CONSEQUENTIAL DAMAGES, ARISING OUT OF THE
 * USE OF THIS CODE.
 *********************************************************************/

typedef struct {   // unpacked structure
  int  i_data;
  real r_data;
} data_t;

module buffer (input  data_t  in,
               output data_t  out);
  //...
endmodule

module chip (/*...*/);

  data_t dint;        // unpacked structure

  struct {            // unpacked structure
    int  i_data;
    real r_data;
  } dout;

  buffer i1 (.in(din),    // legal connection (same typedef type)
             .out(dout)   // illegal connection (not same typedef type)
            );
  //...
endmodule

module test;
  initial begin
    $display("\nExpect error on second port of instance i1 of buffer");
    $display("No simulation results--just checking compilation/elaboration\n");
    $finish;
  end
endmodule
