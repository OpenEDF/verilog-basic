package router_stimulus_pkg;

import uvm_pkg::*;

`include "packet.sv"
`include "packet_da_3.sv"
`include "packet_sequence.sv"

`include "reset_tr.sv"
`include "reset_sequence.sv"

`include "router_input_port_reset_sequence.sv"

endpackage
