module example (/*AUTOARG*/);
   input i;
   output o;

   /*AUTOINPUT*/
   /*AUTOOUTPUT*/
   /*AUTOREG*/
   always @ (/*AUTOSENSE*/) begin
      o = i;
   end

endmodule // example
