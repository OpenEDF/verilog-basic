// # 1. Verilog File Header:


// # 2. Verilog Code style:
module [module_name] (
    [mode] [data_type] [port_names],
    [mode] [data_type] [port_names],
    [mode] [data_type] [port_names]
);



endmodule

// #3. File comment

//--------------------------------------------------------------------------
//
//--------------------------------------------------------------------------
