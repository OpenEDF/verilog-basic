// test bench
`timescale 1ns/1ps
module top_tb();

/* instant pc */
/* instant ram */
/* instant if_id */

/* dispaly mem */

/* clk */


endmodule
