/**********************************************************************
 * while loops
 *
 * Author: Stuart Sutherland
 *
 * (c) Copyright 2003, Sutherland HDL, Inc. *** ALL RIGHTS RESERVED ***
 * www.sutherland-hdl.com
 *
 * Used with permission in the book, "SystemVerilog for Design"
 *  By Stuart Sutherland, Simon Davidmann, and Peter Flake.
 *  Book copyright: 2003, Kluwer Academic Publishers, Norwell, MA, USA
 *  www.wkap.il, ISBN: 0-4020-7530-8
 *
 * Revision History:
 *   1.00 15 Dec 2003 -- original code, as included in book
 *   1.01 10 Jul 2004 -- cleaned up comments, added expected results
 *                       to output messages
 *
 * Caveat: Expected results displayed for this code example are based
 * on an interpretation of the SystemVerilog 3.1 standard by the code
 * author or authors.  At the time of writing, official SystemVerilog
 * validation suites were not available to validate the example.
 *
 * RIGHT TO USE: This code example, or any portion thereof, may be
 * used and distributed without restriction, provided that this entire
 * comment block is included with the example.
 *
 * DISCLAIMER: THIS CODE EXAMPLE IS PROVIDED "AS IS" WITHOUT WARRANTY
 * OF ANY KIND, EITHER EXPRESS OR IMPLIED, INCLUDING, BUT NOT LIMITED
 * TO WARRANTIES OF MERCHANTABILITY, FITNESS OR CORRECTNESS. IN NO
 * EVENT SHALL THE AUTHOR OR AUTHORS BE LIABLE FOR ANY DAMAGES,
 * INCLUDING INCIDENTAL OR CONSEQUENTIAL DAMAGES, ARISING OUT OF THE
 * USE OF THIS CODE.
 *********************************************************************/

module test;
  bit done, OutOfBound;
  bit [11:0] addr;
  bit [15:0] out;
  bit [15:0] mem [0:511];

  always_comb begin
    if (addr < 128 || addr > 255) begin
      done = 0;
      OutOfBound = 1;
      out = mem[128];
      $display("  addr=%0d  done=%b  OutOfBound=%b", addr, done, OutOfBound);
    end
    else while (addr >= 128 && addr <= 255) begin
      if  (addr == 128) begin
        done = 1;
        OutOfBound = 0;
      end
      else begin
        done = 0;
        OutOfBound = 0;
      end
      $display("  addr=%0d  done=%b  OutOfBound=%b", addr, done, OutOfBound);
      out = mem[addr];
      addr -= 1;
    end
  end

  initial begin
    #1 $display("\nSetting addr=5; expect done=0, OutOfBound=1");
       addr = 5;
    #1 $display("\nSetting addr=128; expect done=1, OutOfBound=0");
       addr = 128;
    #1 $display("\nSetting addr=132; expect addr to decrement to 128");
       addr = 132;
    #1 $display("\nSetting addr=300; expect done=0, OutOfBound=1");
       addr = 300;
    #1 $display("");
    $finish;
  end
endmodule
