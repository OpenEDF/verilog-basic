/* what is class in systemverilog and how to use? */

/* define class */

/* object class instance */

/* declare and create */

/* init */



