//--------------------------------------------------------------------------
//                            UVM Lab
//                         openedf.com
//                     Copyright 2023-2024
//
//                     makermuyi@gmail.com
//
//                       License: BSD
//--------------------------------------------------------------------------
//
// Copyright (c) 2020-2021, openedf.com
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS
// "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT
// LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR
// A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE AUTHOR BE
// LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
// SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR
// BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF
// LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF
// THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF
// SUCH DAMAGE.

//--------------------------------------------------------------------------
// Designer: macro
// Brief: The test is at the top of the hierarchical component that initiates
//        the environment component construction
// Change Log:
//--------------------------------------------------------------------------
`ifndef _AHB_LITE_VSEQ_TEST_SV_
`define _AHB_LITE_VSEQ_TEST_SV_

//--------------------------------------------------------------------------
// Include File
//--------------------------------------------------------------------------
`include "ahb_type.svh"
//--------------------------------------------------------------------------
// Class
//--------------------------------------------------------------------------
bit status;
class ahb_lite_vseq_test extends ahb_lite_base_test;

//--------------------------------------------------------------------------
// Design: declare and register
//--------------------------------------------------------------------------
// ahb_lite_system_config sys_cfg;
`uvm_component_utils(ahb_lite_vseq_test)

//--------------------------------------------------------------------------
// Design: declare method
//--------------------------------------------------------------------------
extern function new(string name = "ahb_lite_vseq_test", uvm_component parent = null);
extern virtual task run_phase(uvm_phase phase);

endclass: ahb_lite_vseq_test
//--------------------------------------------------------------------------
// Design: new
//--------------------------------------------------------------------------
function ahb_lite_vseq_test::new(string name = "ahb_lite_vseq_test", uvm_component parent = null);
    super.new(name, parent);
endfunction

//--------------------------------------------------------------------------
// Design: Test DUT
//--------------------------------------------------------------------------
task ahb_lite_vseq_test::run_phase(uvm_phase phase);
    ahb_mst_vseq vseq = ahb_mst_vseq::type_id::create("vseq");

    `uvm_info(get_type_name(), "run phase Entered ...", UVM_HIGH);

    vseq.set_starting_phase(phase);
    vseq.set_automatic_phase_objection(1);

    status = vseq.get_automatic_phase_objection();
    `uvm_info(get_name(), $sformatf("during seq is running, get_automatic_phase_objection: %b", status), UVM_LOW)

    init_seq(vseq);
    vseq.start(null);

    phase.phase_done.set_drain_time(this, 100);
    /* The drop is expected to be matched with an earlier raise */
    `uvm_info(get_type_name(), "run phase Exited ...", UVM_HIGH);
endtask

`endif /* _AHB_LITE_VSEQ_TEST_SV_ */
//--------------------------------------------------------------------------
