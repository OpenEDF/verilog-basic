package test_base_pkg;
import uvm_pkg::*;

`include "packet.sv"
`include "driver.sv"
`include "input_agent.sv"
`include "router_env.sv"
`include "test_base.sv"

endpackage
