//--------------------------------------------------------------------------
//                            UVM Lab
//                         openedf.com
//                     Copyright 2023-2024
//
//                     makermuyi@gmail.com
//
//                       License: BSD
//--------------------------------------------------------------------------
//
// Copyright (c) 2020-2021, openedf.com
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS
// "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT
// LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR
// A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE AUTHOR BE
// LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
// SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR
// BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF
// LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF
// THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF
// SUCH DAMAGE.

//--------------------------------------------------------------------------
// Designer: macro
// Brief: The test is at the top of the hierarchical component that initiates
//        the environment component construction
// Change Log:
//--------------------------------------------------------------------------
`ifndef _AHB_LITE_PIPELINE_TEST_SV_
`define _AHB_LITE_PIPELINE_TEST_SV_

//--------------------------------------------------------------------------
// Include File
//--------------------------------------------------------------------------
`include "ahb_type.svh"
//--------------------------------------------------------------------------
// Class
//--------------------------------------------------------------------------
class ahb_lite_pipeline_test extends ahb_lite_base_test;

//--------------------------------------------------------------------------
// Design: declare and register
//--------------------------------------------------------------------------
ahb_mst_base_seq  mst_seq;
program_ctrl_reg_seq config_seq;
`uvm_component_utils(ahb_lite_pipeline_test)

//--------------------------------------------------------------------------
// Design: declare method
//--------------------------------------------------------------------------
extern function new(string name = "ahb_lite_pipeline_test", uvm_component parent = null);
extern function void build_phase(uvm_phase phase);
extern task configure_phase(uvm_phase phase);
extern task main_phase(uvm_phase phase);

endclass: ahb_lite_pipeline_test
//--------------------------------------------------------------------------
// Design: new
//--------------------------------------------------------------------------
function ahb_lite_pipeline_test::new(string name = "ahb_lite_pipeline_test", uvm_component parent = null);
    super.new(name, parent);
endfunction

//--------------------------------------------------------------------------
// Design: build phase: create and configure of testbench structure
//--------------------------------------------------------------------------
function void ahb_lite_pipeline_test::build_phase(uvm_phase phase);
    `uvm_info(get_type_name(), "IN build_phase...", UVM_HIGH);
    super.build_phase(phase);
    mst_seq = ahb_mst_base_seq::type_id::create("mst_seq");
    config_seq = program_ctrl_reg_seq::type_id::create("config_seq");
endfunction

//--------------------------------------------------------------------------
// Design: Configure the DUT
//--------------------------------------------------------------------------
task ahb_lite_pipeline_test::configure_phase(uvm_phase phase);
    `uvm_info(get_type_name(), " configure_phase Entered...", UVM_HIGH);

    phase.raise_objection(this);
    config_seq.start(ahb_env.mst_agt.mst_seqr);
    phase.drop_objection(this);

    `uvm_info(get_type_name(), "configure_phase Exited...", UVM_HIGH);
endtask

//--------------------------------------------------------------------------
// Design: main phase: stmulate the DUT
//--------------------------------------------------------------------------
task ahb_lite_pipeline_test::main_phase(uvm_phase phase);
    `uvm_info(get_type_name(), "main_phase Entered...", UVM_HIGH);
    phase.raise_objection(this);

    /* Executes this sequence, returning when the sequence has completed  */
    /* main sequence */
    mst_seq.start(ahb_env.mst_agt.mst_seqr);

    /* The drop is expected to be matched with an earlier raise */
    phase.drop_objection(this);
    `uvm_info(get_type_name(), "main_phase Exited...", UVM_HIGH);
endtask

`endif /*_AHB_LITE_PIPELINE_TEST_SV_ */
//--------------------------------------------------------------------------
