/* Arithmetic Operators */

module arithmetic_operators();

initial begin
    $display("5 + 10 = %d", 5 + 10);
    $finish;
end

endmodule
