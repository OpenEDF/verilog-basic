//--------------------------------------------------------------------------
//                         RISC-V Core
//                            V1.0.0
//                         openedf.com
//                     Copyright 2023-2024
//
//                     makermuyi@gmail.com
//
//                       License: BSD
//--------------------------------------------------------------------------
//
// Copyright (c) 2020-2021, openedf.com
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS
// "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT
// LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR
// A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE AUTHOR BE
// LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
// SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR
// BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF
// LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF
// THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF
// SUCH DAMAGE.

//--------------------------------------------------------------------------
// Designer: macro
// Brief: randomination
// Change Log:
//--------------------------------------------------------------------------

//--------------------------------------------------------------------------
// Include File
//--------------------------------------------------------------------------
`include "packet.sv"

//--------------------------------------------------------------------------
// Module
//--------------------------------------------------------------------------
module testebench;
//--------------------------------------------------------------------------
// Ports
//--------------------------------------------------------------------------

//--------------------------------------------------------------------------
// Design: initial and create 
//--------------------------------------------------------------------------
initial begin
    packet pkt;
    pkt = new();
    pkt.addr_range = "small";

    $display("time: %0t constraint_mode = %0d", $time, pkt.address_range.constraint_mode());
    repeat(10) begin
        pkt.randomize();
        $display("time: %0t %s pkt.addr = %0d", $time, pkt.addr_range, pkt.addr);
    end

   $display("-----------------------------------------");
    pkt.address_range.constraint_mode(0);
        $display("time: %0t constraint_mode = %0d", $time, pkt.address_range.constraint_mode());
    pkt.addr_range = "big";
    repeat(10) begin
        pkt.randomize();
        $display("time: %0t %s pkt.addr = %0d", $time, pkt.addr_range, pkt.addr);
    end

   $display("-----------------------------------------");
    pkt.address_range.constraint_mode(1);
        $display("time: %0t constraint_mode = %0d", $time, pkt.address_range.constraint_mode());
    pkt.addr_range = "big";
    repeat(10) begin
        pkt.randomize();
        $display("time: %0t %s pkt.addr = %0d", $time, pkt.addr_range, pkt.addr);
    end
end

endmodule
//--------------------------------------------------------------------------
