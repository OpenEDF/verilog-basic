//--------------------------------------------------------------------------
//                            UVM Lab
//                         openedf.com
//                     Copyright 2023-2024
//
//                     makermuyi@gmail.com
//
//                       License: BSD
//--------------------------------------------------------------------------
//
// Copyright (c) 2020-2021, openedf.com
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS
// "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT
// LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR
// A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE AUTHOR BE
// LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
// SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR
// BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF
// LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF
// THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF
// SUCH DAMAGE.

//--------------------------------------------------------------------------
// Designer: macro
// Brief: interface connection DUT and driver between
// Change Log:
//--------------------------------------------------------------------------

//--------------------------------------------------------------------------
// Include File
//--------------------------------------------------------------------------

//--------------------------------------------------------------------------
// Interface
//--------------------------------------------------------------------------
interface dma_if (
//--------------------------------------------------------------------------
// Port
//--------------------------------------------------------------------------
    input logic clk,
    input logic rst_n
);

//--------------------------------------------------------------------------
// Design: interface signal
//--------------------------------------------------------------------------
logic [31:0] addr;
logic        wr_en;
logic        valid;
logic [31:0] wdata;
logic [31:0] rdata;

//--------------------------------------------------------------------------
// Design: driver interface clocking block
//--------------------------------------------------------------------------
clocking driver_cb @(posedge clk);
    default input #1 output #1;
    output addr;
    output wr_en;
    output valid;
    output wdata;
    input  rdata;
endclocking

//--------------------------------------------------------------------------
// Design: monitor interface clocking block
//--------------------------------------------------------------------------
clocking monitor_cb @(posedge clk);
   default input #1 output #1;
   input addr;
   input wr_en;
   input valid;
   input wdata;
   input rdata;
endclocking

//--------------------------------------------------------------------------
// Design: driver modport
//--------------------------------------------------------------------------
modport DRIVER (clocking driver_cb, input clk, rst_n);

//--------------------------------------------------------------------------
// Design: monitor modport
//--------------------------------------------------------------------------
modport MONITOR (clocking monitor_cb, input clk, rst_n);

endinterface
//--------------------------------------------------------------------------
