//
// Verilog description for cell my_chip, 
// 02/08/14 01:18:08
//
// Precision RTL Synthesis, 2013a.9//


module my_chip ( clk, in, out ) ;

    input clk ;
    input [581:0]in ;
    output [511:0]out ;

    wire [511:0]out_dup_0;
    wire clk_int;
    wire [581:70]in_int;



    OBUF \out_obuf(0)  (.O (out[0]), .I (out_dup_0[0])) ;
    OBUF \out_obuf(1)  (.O (out[1]), .I (out_dup_0[1])) ;
    OBUF \out_obuf(2)  (.O (out[2]), .I (out_dup_0[2])) ;
    OBUF \out_obuf(3)  (.O (out[3]), .I (out_dup_0[3])) ;
    OBUF \out_obuf(4)  (.O (out[4]), .I (out_dup_0[4])) ;
    OBUF \out_obuf(5)  (.O (out[5]), .I (out_dup_0[5])) ;
    OBUF \out_obuf(6)  (.O (out[6]), .I (out_dup_0[6])) ;
    OBUF \out_obuf(7)  (.O (out[7]), .I (out_dup_0[7])) ;
    OBUF \out_obuf(8)  (.O (out[8]), .I (out_dup_0[8])) ;
    OBUF \out_obuf(9)  (.O (out[9]), .I (out_dup_0[9])) ;
    OBUF \out_obuf(10)  (.O (out[10]), .I (out_dup_0[10])) ;
    OBUF \out_obuf(11)  (.O (out[11]), .I (out_dup_0[11])) ;
    OBUF \out_obuf(12)  (.O (out[12]), .I (out_dup_0[12])) ;
    OBUF \out_obuf(13)  (.O (out[13]), .I (out_dup_0[13])) ;
    OBUF \out_obuf(14)  (.O (out[14]), .I (out_dup_0[14])) ;
    OBUF \out_obuf(15)  (.O (out[15]), .I (out_dup_0[15])) ;
    OBUF \out_obuf(16)  (.O (out[16]), .I (out_dup_0[16])) ;
    OBUF \out_obuf(17)  (.O (out[17]), .I (out_dup_0[17])) ;
    OBUF \out_obuf(18)  (.O (out[18]), .I (out_dup_0[18])) ;
    OBUF \out_obuf(19)  (.O (out[19]), .I (out_dup_0[19])) ;
    OBUF \out_obuf(20)  (.O (out[20]), .I (out_dup_0[20])) ;
    OBUF \out_obuf(21)  (.O (out[21]), .I (out_dup_0[21])) ;
    OBUF \out_obuf(22)  (.O (out[22]), .I (out_dup_0[22])) ;
    OBUF \out_obuf(23)  (.O (out[23]), .I (out_dup_0[23])) ;
    OBUF \out_obuf(24)  (.O (out[24]), .I (out_dup_0[24])) ;
    OBUF \out_obuf(25)  (.O (out[25]), .I (out_dup_0[25])) ;
    OBUF \out_obuf(26)  (.O (out[26]), .I (out_dup_0[26])) ;
    OBUF \out_obuf(27)  (.O (out[27]), .I (out_dup_0[27])) ;
    OBUF \out_obuf(28)  (.O (out[28]), .I (out_dup_0[28])) ;
    OBUF \out_obuf(29)  (.O (out[29]), .I (out_dup_0[29])) ;
    OBUF \out_obuf(30)  (.O (out[30]), .I (out_dup_0[30])) ;
    OBUF \out_obuf(31)  (.O (out[31]), .I (out_dup_0[31])) ;
    OBUF \out_obuf(32)  (.O (out[32]), .I (out_dup_0[32])) ;
    OBUF \out_obuf(33)  (.O (out[33]), .I (out_dup_0[33])) ;
    OBUF \out_obuf(34)  (.O (out[34]), .I (out_dup_0[34])) ;
    OBUF \out_obuf(35)  (.O (out[35]), .I (out_dup_0[35])) ;
    OBUF \out_obuf(36)  (.O (out[36]), .I (out_dup_0[36])) ;
    OBUF \out_obuf(37)  (.O (out[37]), .I (out_dup_0[37])) ;
    OBUF \out_obuf(38)  (.O (out[38]), .I (out_dup_0[38])) ;
    OBUF \out_obuf(39)  (.O (out[39]), .I (out_dup_0[39])) ;
    OBUF \out_obuf(40)  (.O (out[40]), .I (out_dup_0[40])) ;
    OBUF \out_obuf(41)  (.O (out[41]), .I (out_dup_0[41])) ;
    OBUF \out_obuf(42)  (.O (out[42]), .I (out_dup_0[42])) ;
    OBUF \out_obuf(43)  (.O (out[43]), .I (out_dup_0[43])) ;
    OBUF \out_obuf(44)  (.O (out[44]), .I (out_dup_0[44])) ;
    OBUF \out_obuf(45)  (.O (out[45]), .I (out_dup_0[45])) ;
    OBUF \out_obuf(46)  (.O (out[46]), .I (out_dup_0[46])) ;
    OBUF \out_obuf(47)  (.O (out[47]), .I (out_dup_0[47])) ;
    OBUF \out_obuf(48)  (.O (out[48]), .I (out_dup_0[48])) ;
    OBUF \out_obuf(49)  (.O (out[49]), .I (out_dup_0[49])) ;
    OBUF \out_obuf(50)  (.O (out[50]), .I (out_dup_0[50])) ;
    OBUF \out_obuf(51)  (.O (out[51]), .I (out_dup_0[51])) ;
    OBUF \out_obuf(52)  (.O (out[52]), .I (out_dup_0[52])) ;
    OBUF \out_obuf(53)  (.O (out[53]), .I (out_dup_0[53])) ;
    OBUF \out_obuf(54)  (.O (out[54]), .I (out_dup_0[54])) ;
    OBUF \out_obuf(55)  (.O (out[55]), .I (out_dup_0[55])) ;
    OBUF \out_obuf(56)  (.O (out[56]), .I (out_dup_0[56])) ;
    OBUF \out_obuf(57)  (.O (out[57]), .I (out_dup_0[57])) ;
    OBUF \out_obuf(58)  (.O (out[58]), .I (out_dup_0[58])) ;
    OBUF \out_obuf(59)  (.O (out[59]), .I (out_dup_0[59])) ;
    OBUF \out_obuf(60)  (.O (out[60]), .I (out_dup_0[60])) ;
    OBUF \out_obuf(61)  (.O (out[61]), .I (out_dup_0[61])) ;
    OBUF \out_obuf(62)  (.O (out[62]), .I (out_dup_0[62])) ;
    OBUF \out_obuf(63)  (.O (out[63]), .I (out_dup_0[63])) ;
    OBUF \out_obuf(64)  (.O (out[64]), .I (out_dup_0[64])) ;
    OBUF \out_obuf(65)  (.O (out[65]), .I (out_dup_0[65])) ;
    OBUF \out_obuf(66)  (.O (out[66]), .I (out_dup_0[66])) ;
    OBUF \out_obuf(67)  (.O (out[67]), .I (out_dup_0[67])) ;
    OBUF \out_obuf(68)  (.O (out[68]), .I (out_dup_0[68])) ;
    OBUF \out_obuf(69)  (.O (out[69]), .I (out_dup_0[69])) ;
    OBUF \out_obuf(70)  (.O (out[70]), .I (out_dup_0[70])) ;
    OBUF \out_obuf(71)  (.O (out[71]), .I (out_dup_0[71])) ;
    OBUF \out_obuf(72)  (.O (out[72]), .I (out_dup_0[72])) ;
    OBUF \out_obuf(73)  (.O (out[73]), .I (out_dup_0[73])) ;
    OBUF \out_obuf(74)  (.O (out[74]), .I (out_dup_0[74])) ;
    OBUF \out_obuf(75)  (.O (out[75]), .I (out_dup_0[75])) ;
    OBUF \out_obuf(76)  (.O (out[76]), .I (out_dup_0[76])) ;
    OBUF \out_obuf(77)  (.O (out[77]), .I (out_dup_0[77])) ;
    OBUF \out_obuf(78)  (.O (out[78]), .I (out_dup_0[78])) ;
    OBUF \out_obuf(79)  (.O (out[79]), .I (out_dup_0[79])) ;
    OBUF \out_obuf(80)  (.O (out[80]), .I (out_dup_0[80])) ;
    OBUF \out_obuf(81)  (.O (out[81]), .I (out_dup_0[81])) ;
    OBUF \out_obuf(82)  (.O (out[82]), .I (out_dup_0[82])) ;
    OBUF \out_obuf(83)  (.O (out[83]), .I (out_dup_0[83])) ;
    OBUF \out_obuf(84)  (.O (out[84]), .I (out_dup_0[84])) ;
    OBUF \out_obuf(85)  (.O (out[85]), .I (out_dup_0[85])) ;
    OBUF \out_obuf(86)  (.O (out[86]), .I (out_dup_0[86])) ;
    OBUF \out_obuf(87)  (.O (out[87]), .I (out_dup_0[87])) ;
    OBUF \out_obuf(88)  (.O (out[88]), .I (out_dup_0[88])) ;
    OBUF \out_obuf(89)  (.O (out[89]), .I (out_dup_0[89])) ;
    OBUF \out_obuf(90)  (.O (out[90]), .I (out_dup_0[90])) ;
    OBUF \out_obuf(91)  (.O (out[91]), .I (out_dup_0[91])) ;
    OBUF \out_obuf(92)  (.O (out[92]), .I (out_dup_0[92])) ;
    OBUF \out_obuf(93)  (.O (out[93]), .I (out_dup_0[93])) ;
    OBUF \out_obuf(94)  (.O (out[94]), .I (out_dup_0[94])) ;
    OBUF \out_obuf(95)  (.O (out[95]), .I (out_dup_0[95])) ;
    OBUF \out_obuf(96)  (.O (out[96]), .I (out_dup_0[96])) ;
    OBUF \out_obuf(97)  (.O (out[97]), .I (out_dup_0[97])) ;
    OBUF \out_obuf(98)  (.O (out[98]), .I (out_dup_0[98])) ;
    OBUF \out_obuf(99)  (.O (out[99]), .I (out_dup_0[99])) ;
    OBUF \out_obuf(100)  (.O (out[100]), .I (out_dup_0[100])) ;
    OBUF \out_obuf(101)  (.O (out[101]), .I (out_dup_0[101])) ;
    OBUF \out_obuf(102)  (.O (out[102]), .I (out_dup_0[102])) ;
    OBUF \out_obuf(103)  (.O (out[103]), .I (out_dup_0[103])) ;
    OBUF \out_obuf(104)  (.O (out[104]), .I (out_dup_0[104])) ;
    OBUF \out_obuf(105)  (.O (out[105]), .I (out_dup_0[105])) ;
    OBUF \out_obuf(106)  (.O (out[106]), .I (out_dup_0[106])) ;
    OBUF \out_obuf(107)  (.O (out[107]), .I (out_dup_0[107])) ;
    OBUF \out_obuf(108)  (.O (out[108]), .I (out_dup_0[108])) ;
    OBUF \out_obuf(109)  (.O (out[109]), .I (out_dup_0[109])) ;
    OBUF \out_obuf(110)  (.O (out[110]), .I (out_dup_0[110])) ;
    OBUF \out_obuf(111)  (.O (out[111]), .I (out_dup_0[111])) ;
    OBUF \out_obuf(112)  (.O (out[112]), .I (out_dup_0[112])) ;
    OBUF \out_obuf(113)  (.O (out[113]), .I (out_dup_0[113])) ;
    OBUF \out_obuf(114)  (.O (out[114]), .I (out_dup_0[114])) ;
    OBUF \out_obuf(115)  (.O (out[115]), .I (out_dup_0[115])) ;
    OBUF \out_obuf(116)  (.O (out[116]), .I (out_dup_0[116])) ;
    OBUF \out_obuf(117)  (.O (out[117]), .I (out_dup_0[117])) ;
    OBUF \out_obuf(118)  (.O (out[118]), .I (out_dup_0[118])) ;
    OBUF \out_obuf(119)  (.O (out[119]), .I (out_dup_0[119])) ;
    OBUF \out_obuf(120)  (.O (out[120]), .I (out_dup_0[120])) ;
    OBUF \out_obuf(121)  (.O (out[121]), .I (out_dup_0[121])) ;
    OBUF \out_obuf(122)  (.O (out[122]), .I (out_dup_0[122])) ;
    OBUF \out_obuf(123)  (.O (out[123]), .I (out_dup_0[123])) ;
    OBUF \out_obuf(124)  (.O (out[124]), .I (out_dup_0[124])) ;
    OBUF \out_obuf(125)  (.O (out[125]), .I (out_dup_0[125])) ;
    OBUF \out_obuf(126)  (.O (out[126]), .I (out_dup_0[126])) ;
    OBUF \out_obuf(127)  (.O (out[127]), .I (out_dup_0[127])) ;
    OBUF \out_obuf(128)  (.O (out[128]), .I (out_dup_0[128])) ;
    OBUF \out_obuf(129)  (.O (out[129]), .I (out_dup_0[129])) ;
    OBUF \out_obuf(130)  (.O (out[130]), .I (out_dup_0[130])) ;
    OBUF \out_obuf(131)  (.O (out[131]), .I (out_dup_0[131])) ;
    OBUF \out_obuf(132)  (.O (out[132]), .I (out_dup_0[132])) ;
    OBUF \out_obuf(133)  (.O (out[133]), .I (out_dup_0[133])) ;
    OBUF \out_obuf(134)  (.O (out[134]), .I (out_dup_0[134])) ;
    OBUF \out_obuf(135)  (.O (out[135]), .I (out_dup_0[135])) ;
    OBUF \out_obuf(136)  (.O (out[136]), .I (out_dup_0[136])) ;
    OBUF \out_obuf(137)  (.O (out[137]), .I (out_dup_0[137])) ;
    OBUF \out_obuf(138)  (.O (out[138]), .I (out_dup_0[138])) ;
    OBUF \out_obuf(139)  (.O (out[139]), .I (out_dup_0[139])) ;
    OBUF \out_obuf(140)  (.O (out[140]), .I (out_dup_0[140])) ;
    OBUF \out_obuf(141)  (.O (out[141]), .I (out_dup_0[141])) ;
    OBUF \out_obuf(142)  (.O (out[142]), .I (out_dup_0[142])) ;
    OBUF \out_obuf(143)  (.O (out[143]), .I (out_dup_0[143])) ;
    OBUF \out_obuf(144)  (.O (out[144]), .I (out_dup_0[144])) ;
    OBUF \out_obuf(145)  (.O (out[145]), .I (out_dup_0[145])) ;
    OBUF \out_obuf(146)  (.O (out[146]), .I (out_dup_0[146])) ;
    OBUF \out_obuf(147)  (.O (out[147]), .I (out_dup_0[147])) ;
    OBUF \out_obuf(148)  (.O (out[148]), .I (out_dup_0[148])) ;
    OBUF \out_obuf(149)  (.O (out[149]), .I (out_dup_0[149])) ;
    OBUF \out_obuf(150)  (.O (out[150]), .I (out_dup_0[150])) ;
    OBUF \out_obuf(151)  (.O (out[151]), .I (out_dup_0[151])) ;
    OBUF \out_obuf(152)  (.O (out[152]), .I (out_dup_0[152])) ;
    OBUF \out_obuf(153)  (.O (out[153]), .I (out_dup_0[153])) ;
    OBUF \out_obuf(154)  (.O (out[154]), .I (out_dup_0[154])) ;
    OBUF \out_obuf(155)  (.O (out[155]), .I (out_dup_0[155])) ;
    OBUF \out_obuf(156)  (.O (out[156]), .I (out_dup_0[156])) ;
    OBUF \out_obuf(157)  (.O (out[157]), .I (out_dup_0[157])) ;
    OBUF \out_obuf(158)  (.O (out[158]), .I (out_dup_0[158])) ;
    OBUF \out_obuf(159)  (.O (out[159]), .I (out_dup_0[159])) ;
    OBUF \out_obuf(160)  (.O (out[160]), .I (out_dup_0[160])) ;
    OBUF \out_obuf(161)  (.O (out[161]), .I (out_dup_0[161])) ;
    OBUF \out_obuf(162)  (.O (out[162]), .I (out_dup_0[162])) ;
    OBUF \out_obuf(163)  (.O (out[163]), .I (out_dup_0[163])) ;
    OBUF \out_obuf(164)  (.O (out[164]), .I (out_dup_0[164])) ;
    OBUF \out_obuf(165)  (.O (out[165]), .I (out_dup_0[165])) ;
    OBUF \out_obuf(166)  (.O (out[166]), .I (out_dup_0[166])) ;
    OBUF \out_obuf(167)  (.O (out[167]), .I (out_dup_0[167])) ;
    OBUF \out_obuf(168)  (.O (out[168]), .I (out_dup_0[168])) ;
    OBUF \out_obuf(169)  (.O (out[169]), .I (out_dup_0[169])) ;
    OBUF \out_obuf(170)  (.O (out[170]), .I (out_dup_0[170])) ;
    OBUF \out_obuf(171)  (.O (out[171]), .I (out_dup_0[171])) ;
    OBUF \out_obuf(172)  (.O (out[172]), .I (out_dup_0[172])) ;
    OBUF \out_obuf(173)  (.O (out[173]), .I (out_dup_0[173])) ;
    OBUF \out_obuf(174)  (.O (out[174]), .I (out_dup_0[174])) ;
    OBUF \out_obuf(175)  (.O (out[175]), .I (out_dup_0[175])) ;
    OBUF \out_obuf(176)  (.O (out[176]), .I (out_dup_0[176])) ;
    OBUF \out_obuf(177)  (.O (out[177]), .I (out_dup_0[177])) ;
    OBUF \out_obuf(178)  (.O (out[178]), .I (out_dup_0[178])) ;
    OBUF \out_obuf(179)  (.O (out[179]), .I (out_dup_0[179])) ;
    OBUF \out_obuf(180)  (.O (out[180]), .I (out_dup_0[180])) ;
    OBUF \out_obuf(181)  (.O (out[181]), .I (out_dup_0[181])) ;
    OBUF \out_obuf(182)  (.O (out[182]), .I (out_dup_0[182])) ;
    OBUF \out_obuf(183)  (.O (out[183]), .I (out_dup_0[183])) ;
    OBUF \out_obuf(184)  (.O (out[184]), .I (out_dup_0[184])) ;
    OBUF \out_obuf(185)  (.O (out[185]), .I (out_dup_0[185])) ;
    OBUF \out_obuf(186)  (.O (out[186]), .I (out_dup_0[186])) ;
    OBUF \out_obuf(187)  (.O (out[187]), .I (out_dup_0[187])) ;
    OBUF \out_obuf(188)  (.O (out[188]), .I (out_dup_0[188])) ;
    OBUF \out_obuf(189)  (.O (out[189]), .I (out_dup_0[189])) ;
    OBUF \out_obuf(190)  (.O (out[190]), .I (out_dup_0[190])) ;
    OBUF \out_obuf(191)  (.O (out[191]), .I (out_dup_0[191])) ;
    OBUF \out_obuf(192)  (.O (out[192]), .I (out_dup_0[192])) ;
    OBUF \out_obuf(193)  (.O (out[193]), .I (out_dup_0[193])) ;
    OBUF \out_obuf(194)  (.O (out[194]), .I (out_dup_0[194])) ;
    OBUF \out_obuf(195)  (.O (out[195]), .I (out_dup_0[195])) ;
    OBUF \out_obuf(196)  (.O (out[196]), .I (out_dup_0[196])) ;
    OBUF \out_obuf(197)  (.O (out[197]), .I (out_dup_0[197])) ;
    OBUF \out_obuf(198)  (.O (out[198]), .I (out_dup_0[198])) ;
    OBUF \out_obuf(199)  (.O (out[199]), .I (out_dup_0[199])) ;
    OBUF \out_obuf(200)  (.O (out[200]), .I (out_dup_0[200])) ;
    OBUF \out_obuf(201)  (.O (out[201]), .I (out_dup_0[201])) ;
    OBUF \out_obuf(202)  (.O (out[202]), .I (out_dup_0[202])) ;
    OBUF \out_obuf(203)  (.O (out[203]), .I (out_dup_0[203])) ;
    OBUF \out_obuf(204)  (.O (out[204]), .I (out_dup_0[204])) ;
    OBUF \out_obuf(205)  (.O (out[205]), .I (out_dup_0[205])) ;
    OBUF \out_obuf(206)  (.O (out[206]), .I (out_dup_0[206])) ;
    OBUF \out_obuf(207)  (.O (out[207]), .I (out_dup_0[207])) ;
    OBUF \out_obuf(208)  (.O (out[208]), .I (out_dup_0[208])) ;
    OBUF \out_obuf(209)  (.O (out[209]), .I (out_dup_0[209])) ;
    OBUF \out_obuf(210)  (.O (out[210]), .I (out_dup_0[210])) ;
    OBUF \out_obuf(211)  (.O (out[211]), .I (out_dup_0[211])) ;
    OBUF \out_obuf(212)  (.O (out[212]), .I (out_dup_0[212])) ;
    OBUF \out_obuf(213)  (.O (out[213]), .I (out_dup_0[213])) ;
    OBUF \out_obuf(214)  (.O (out[214]), .I (out_dup_0[214])) ;
    OBUF \out_obuf(215)  (.O (out[215]), .I (out_dup_0[215])) ;
    OBUF \out_obuf(216)  (.O (out[216]), .I (out_dup_0[216])) ;
    OBUF \out_obuf(217)  (.O (out[217]), .I (out_dup_0[217])) ;
    OBUF \out_obuf(218)  (.O (out[218]), .I (out_dup_0[218])) ;
    OBUF \out_obuf(219)  (.O (out[219]), .I (out_dup_0[219])) ;
    OBUF \out_obuf(220)  (.O (out[220]), .I (out_dup_0[220])) ;
    OBUF \out_obuf(221)  (.O (out[221]), .I (out_dup_0[221])) ;
    OBUF \out_obuf(222)  (.O (out[222]), .I (out_dup_0[222])) ;
    OBUF \out_obuf(223)  (.O (out[223]), .I (out_dup_0[223])) ;
    OBUF \out_obuf(224)  (.O (out[224]), .I (out_dup_0[224])) ;
    OBUF \out_obuf(225)  (.O (out[225]), .I (out_dup_0[225])) ;
    OBUF \out_obuf(226)  (.O (out[226]), .I (out_dup_0[226])) ;
    OBUF \out_obuf(227)  (.O (out[227]), .I (out_dup_0[227])) ;
    OBUF \out_obuf(228)  (.O (out[228]), .I (out_dup_0[228])) ;
    OBUF \out_obuf(229)  (.O (out[229]), .I (out_dup_0[229])) ;
    OBUF \out_obuf(230)  (.O (out[230]), .I (out_dup_0[230])) ;
    OBUF \out_obuf(231)  (.O (out[231]), .I (out_dup_0[231])) ;
    OBUF \out_obuf(232)  (.O (out[232]), .I (out_dup_0[232])) ;
    OBUF \out_obuf(233)  (.O (out[233]), .I (out_dup_0[233])) ;
    OBUF \out_obuf(234)  (.O (out[234]), .I (out_dup_0[234])) ;
    OBUF \out_obuf(235)  (.O (out[235]), .I (out_dup_0[235])) ;
    OBUF \out_obuf(236)  (.O (out[236]), .I (out_dup_0[236])) ;
    OBUF \out_obuf(237)  (.O (out[237]), .I (out_dup_0[237])) ;
    OBUF \out_obuf(238)  (.O (out[238]), .I (out_dup_0[238])) ;
    OBUF \out_obuf(239)  (.O (out[239]), .I (out_dup_0[239])) ;
    OBUF \out_obuf(240)  (.O (out[240]), .I (out_dup_0[240])) ;
    OBUF \out_obuf(241)  (.O (out[241]), .I (out_dup_0[241])) ;
    OBUF \out_obuf(242)  (.O (out[242]), .I (out_dup_0[242])) ;
    OBUF \out_obuf(243)  (.O (out[243]), .I (out_dup_0[243])) ;
    OBUF \out_obuf(244)  (.O (out[244]), .I (out_dup_0[244])) ;
    OBUF \out_obuf(245)  (.O (out[245]), .I (out_dup_0[245])) ;
    OBUF \out_obuf(246)  (.O (out[246]), .I (out_dup_0[246])) ;
    OBUF \out_obuf(247)  (.O (out[247]), .I (out_dup_0[247])) ;
    OBUF \out_obuf(248)  (.O (out[248]), .I (out_dup_0[248])) ;
    OBUF \out_obuf(249)  (.O (out[249]), .I (out_dup_0[249])) ;
    OBUF \out_obuf(250)  (.O (out[250]), .I (out_dup_0[250])) ;
    OBUF \out_obuf(251)  (.O (out[251]), .I (out_dup_0[251])) ;
    OBUF \out_obuf(252)  (.O (out[252]), .I (out_dup_0[252])) ;
    OBUF \out_obuf(253)  (.O (out[253]), .I (out_dup_0[253])) ;
    OBUF \out_obuf(254)  (.O (out[254]), .I (out_dup_0[254])) ;
    OBUF \out_obuf(255)  (.O (out[255]), .I (out_dup_0[255])) ;
    OBUF \out_obuf(256)  (.O (out[256]), .I (out_dup_0[256])) ;
    OBUF \out_obuf(257)  (.O (out[257]), .I (out_dup_0[257])) ;
    OBUF \out_obuf(258)  (.O (out[258]), .I (out_dup_0[258])) ;
    OBUF \out_obuf(259)  (.O (out[259]), .I (out_dup_0[259])) ;
    OBUF \out_obuf(260)  (.O (out[260]), .I (out_dup_0[260])) ;
    OBUF \out_obuf(261)  (.O (out[261]), .I (out_dup_0[261])) ;
    OBUF \out_obuf(262)  (.O (out[262]), .I (out_dup_0[262])) ;
    OBUF \out_obuf(263)  (.O (out[263]), .I (out_dup_0[263])) ;
    OBUF \out_obuf(264)  (.O (out[264]), .I (out_dup_0[264])) ;
    OBUF \out_obuf(265)  (.O (out[265]), .I (out_dup_0[265])) ;
    OBUF \out_obuf(266)  (.O (out[266]), .I (out_dup_0[266])) ;
    OBUF \out_obuf(267)  (.O (out[267]), .I (out_dup_0[267])) ;
    OBUF \out_obuf(268)  (.O (out[268]), .I (out_dup_0[268])) ;
    OBUF \out_obuf(269)  (.O (out[269]), .I (out_dup_0[269])) ;
    OBUF \out_obuf(270)  (.O (out[270]), .I (out_dup_0[270])) ;
    OBUF \out_obuf(271)  (.O (out[271]), .I (out_dup_0[271])) ;
    OBUF \out_obuf(272)  (.O (out[272]), .I (out_dup_0[272])) ;
    OBUF \out_obuf(273)  (.O (out[273]), .I (out_dup_0[273])) ;
    OBUF \out_obuf(274)  (.O (out[274]), .I (out_dup_0[274])) ;
    OBUF \out_obuf(275)  (.O (out[275]), .I (out_dup_0[275])) ;
    OBUF \out_obuf(276)  (.O (out[276]), .I (out_dup_0[276])) ;
    OBUF \out_obuf(277)  (.O (out[277]), .I (out_dup_0[277])) ;
    OBUF \out_obuf(278)  (.O (out[278]), .I (out_dup_0[278])) ;
    OBUF \out_obuf(279)  (.O (out[279]), .I (out_dup_0[279])) ;
    OBUF \out_obuf(280)  (.O (out[280]), .I (out_dup_0[280])) ;
    OBUF \out_obuf(281)  (.O (out[281]), .I (out_dup_0[281])) ;
    OBUF \out_obuf(282)  (.O (out[282]), .I (out_dup_0[282])) ;
    OBUF \out_obuf(283)  (.O (out[283]), .I (out_dup_0[283])) ;
    OBUF \out_obuf(284)  (.O (out[284]), .I (out_dup_0[284])) ;
    OBUF \out_obuf(285)  (.O (out[285]), .I (out_dup_0[285])) ;
    OBUF \out_obuf(286)  (.O (out[286]), .I (out_dup_0[286])) ;
    OBUF \out_obuf(287)  (.O (out[287]), .I (out_dup_0[287])) ;
    OBUF \out_obuf(288)  (.O (out[288]), .I (out_dup_0[288])) ;
    OBUF \out_obuf(289)  (.O (out[289]), .I (out_dup_0[289])) ;
    OBUF \out_obuf(290)  (.O (out[290]), .I (out_dup_0[290])) ;
    OBUF \out_obuf(291)  (.O (out[291]), .I (out_dup_0[291])) ;
    OBUF \out_obuf(292)  (.O (out[292]), .I (out_dup_0[292])) ;
    OBUF \out_obuf(293)  (.O (out[293]), .I (out_dup_0[293])) ;
    OBUF \out_obuf(294)  (.O (out[294]), .I (out_dup_0[294])) ;
    OBUF \out_obuf(295)  (.O (out[295]), .I (out_dup_0[295])) ;
    OBUF \out_obuf(296)  (.O (out[296]), .I (out_dup_0[296])) ;
    OBUF \out_obuf(297)  (.O (out[297]), .I (out_dup_0[297])) ;
    OBUF \out_obuf(298)  (.O (out[298]), .I (out_dup_0[298])) ;
    OBUF \out_obuf(299)  (.O (out[299]), .I (out_dup_0[299])) ;
    OBUF \out_obuf(300)  (.O (out[300]), .I (out_dup_0[300])) ;
    OBUF \out_obuf(301)  (.O (out[301]), .I (out_dup_0[301])) ;
    OBUF \out_obuf(302)  (.O (out[302]), .I (out_dup_0[302])) ;
    OBUF \out_obuf(303)  (.O (out[303]), .I (out_dup_0[303])) ;
    OBUF \out_obuf(304)  (.O (out[304]), .I (out_dup_0[304])) ;
    OBUF \out_obuf(305)  (.O (out[305]), .I (out_dup_0[305])) ;
    OBUF \out_obuf(306)  (.O (out[306]), .I (out_dup_0[306])) ;
    OBUF \out_obuf(307)  (.O (out[307]), .I (out_dup_0[307])) ;
    OBUF \out_obuf(308)  (.O (out[308]), .I (out_dup_0[308])) ;
    OBUF \out_obuf(309)  (.O (out[309]), .I (out_dup_0[309])) ;
    OBUF \out_obuf(310)  (.O (out[310]), .I (out_dup_0[310])) ;
    OBUF \out_obuf(311)  (.O (out[311]), .I (out_dup_0[311])) ;
    OBUF \out_obuf(312)  (.O (out[312]), .I (out_dup_0[312])) ;
    OBUF \out_obuf(313)  (.O (out[313]), .I (out_dup_0[313])) ;
    OBUF \out_obuf(314)  (.O (out[314]), .I (out_dup_0[314])) ;
    OBUF \out_obuf(315)  (.O (out[315]), .I (out_dup_0[315])) ;
    OBUF \out_obuf(316)  (.O (out[316]), .I (out_dup_0[316])) ;
    OBUF \out_obuf(317)  (.O (out[317]), .I (out_dup_0[317])) ;
    OBUF \out_obuf(318)  (.O (out[318]), .I (out_dup_0[318])) ;
    OBUF \out_obuf(319)  (.O (out[319]), .I (out_dup_0[319])) ;
    OBUF \out_obuf(320)  (.O (out[320]), .I (out_dup_0[320])) ;
    OBUF \out_obuf(321)  (.O (out[321]), .I (out_dup_0[321])) ;
    OBUF \out_obuf(322)  (.O (out[322]), .I (out_dup_0[322])) ;
    OBUF \out_obuf(323)  (.O (out[323]), .I (out_dup_0[323])) ;
    OBUF \out_obuf(324)  (.O (out[324]), .I (out_dup_0[324])) ;
    OBUF \out_obuf(325)  (.O (out[325]), .I (out_dup_0[325])) ;
    OBUF \out_obuf(326)  (.O (out[326]), .I (out_dup_0[326])) ;
    OBUF \out_obuf(327)  (.O (out[327]), .I (out_dup_0[327])) ;
    OBUF \out_obuf(328)  (.O (out[328]), .I (out_dup_0[328])) ;
    OBUF \out_obuf(329)  (.O (out[329]), .I (out_dup_0[329])) ;
    OBUF \out_obuf(330)  (.O (out[330]), .I (out_dup_0[330])) ;
    OBUF \out_obuf(331)  (.O (out[331]), .I (out_dup_0[331])) ;
    OBUF \out_obuf(332)  (.O (out[332]), .I (out_dup_0[332])) ;
    OBUF \out_obuf(333)  (.O (out[333]), .I (out_dup_0[333])) ;
    OBUF \out_obuf(334)  (.O (out[334]), .I (out_dup_0[334])) ;
    OBUF \out_obuf(335)  (.O (out[335]), .I (out_dup_0[335])) ;
    OBUF \out_obuf(336)  (.O (out[336]), .I (out_dup_0[336])) ;
    OBUF \out_obuf(337)  (.O (out[337]), .I (out_dup_0[337])) ;
    OBUF \out_obuf(338)  (.O (out[338]), .I (out_dup_0[338])) ;
    OBUF \out_obuf(339)  (.O (out[339]), .I (out_dup_0[339])) ;
    OBUF \out_obuf(340)  (.O (out[340]), .I (out_dup_0[340])) ;
    OBUF \out_obuf(341)  (.O (out[341]), .I (out_dup_0[341])) ;
    OBUF \out_obuf(342)  (.O (out[342]), .I (out_dup_0[342])) ;
    OBUF \out_obuf(343)  (.O (out[343]), .I (out_dup_0[343])) ;
    OBUF \out_obuf(344)  (.O (out[344]), .I (out_dup_0[344])) ;
    OBUF \out_obuf(345)  (.O (out[345]), .I (out_dup_0[345])) ;
    OBUF \out_obuf(346)  (.O (out[346]), .I (out_dup_0[346])) ;
    OBUF \out_obuf(347)  (.O (out[347]), .I (out_dup_0[347])) ;
    OBUF \out_obuf(348)  (.O (out[348]), .I (out_dup_0[348])) ;
    OBUF \out_obuf(349)  (.O (out[349]), .I (out_dup_0[349])) ;
    OBUF \out_obuf(350)  (.O (out[350]), .I (out_dup_0[350])) ;
    OBUF \out_obuf(351)  (.O (out[351]), .I (out_dup_0[351])) ;
    OBUF \out_obuf(352)  (.O (out[352]), .I (out_dup_0[352])) ;
    OBUF \out_obuf(353)  (.O (out[353]), .I (out_dup_0[353])) ;
    OBUF \out_obuf(354)  (.O (out[354]), .I (out_dup_0[354])) ;
    OBUF \out_obuf(355)  (.O (out[355]), .I (out_dup_0[355])) ;
    OBUF \out_obuf(356)  (.O (out[356]), .I (out_dup_0[356])) ;
    OBUF \out_obuf(357)  (.O (out[357]), .I (out_dup_0[357])) ;
    OBUF \out_obuf(358)  (.O (out[358]), .I (out_dup_0[358])) ;
    OBUF \out_obuf(359)  (.O (out[359]), .I (out_dup_0[359])) ;
    OBUF \out_obuf(360)  (.O (out[360]), .I (out_dup_0[360])) ;
    OBUF \out_obuf(361)  (.O (out[361]), .I (out_dup_0[361])) ;
    OBUF \out_obuf(362)  (.O (out[362]), .I (out_dup_0[362])) ;
    OBUF \out_obuf(363)  (.O (out[363]), .I (out_dup_0[363])) ;
    OBUF \out_obuf(364)  (.O (out[364]), .I (out_dup_0[364])) ;
    OBUF \out_obuf(365)  (.O (out[365]), .I (out_dup_0[365])) ;
    OBUF \out_obuf(366)  (.O (out[366]), .I (out_dup_0[366])) ;
    OBUF \out_obuf(367)  (.O (out[367]), .I (out_dup_0[367])) ;
    OBUF \out_obuf(368)  (.O (out[368]), .I (out_dup_0[368])) ;
    OBUF \out_obuf(369)  (.O (out[369]), .I (out_dup_0[369])) ;
    OBUF \out_obuf(370)  (.O (out[370]), .I (out_dup_0[370])) ;
    OBUF \out_obuf(371)  (.O (out[371]), .I (out_dup_0[371])) ;
    OBUF \out_obuf(372)  (.O (out[372]), .I (out_dup_0[372])) ;
    OBUF \out_obuf(373)  (.O (out[373]), .I (out_dup_0[373])) ;
    OBUF \out_obuf(374)  (.O (out[374]), .I (out_dup_0[374])) ;
    OBUF \out_obuf(375)  (.O (out[375]), .I (out_dup_0[375])) ;
    OBUF \out_obuf(376)  (.O (out[376]), .I (out_dup_0[376])) ;
    OBUF \out_obuf(377)  (.O (out[377]), .I (out_dup_0[377])) ;
    OBUF \out_obuf(378)  (.O (out[378]), .I (out_dup_0[378])) ;
    OBUF \out_obuf(379)  (.O (out[379]), .I (out_dup_0[379])) ;
    OBUF \out_obuf(380)  (.O (out[380]), .I (out_dup_0[380])) ;
    OBUF \out_obuf(381)  (.O (out[381]), .I (out_dup_0[381])) ;
    OBUF \out_obuf(382)  (.O (out[382]), .I (out_dup_0[382])) ;
    OBUF \out_obuf(383)  (.O (out[383]), .I (out_dup_0[383])) ;
    OBUF \out_obuf(384)  (.O (out[384]), .I (out_dup_0[384])) ;
    OBUF \out_obuf(385)  (.O (out[385]), .I (out_dup_0[385])) ;
    OBUF \out_obuf(386)  (.O (out[386]), .I (out_dup_0[386])) ;
    OBUF \out_obuf(387)  (.O (out[387]), .I (out_dup_0[387])) ;
    OBUF \out_obuf(388)  (.O (out[388]), .I (out_dup_0[388])) ;
    OBUF \out_obuf(389)  (.O (out[389]), .I (out_dup_0[389])) ;
    OBUF \out_obuf(390)  (.O (out[390]), .I (out_dup_0[390])) ;
    OBUF \out_obuf(391)  (.O (out[391]), .I (out_dup_0[391])) ;
    OBUF \out_obuf(392)  (.O (out[392]), .I (out_dup_0[392])) ;
    OBUF \out_obuf(393)  (.O (out[393]), .I (out_dup_0[393])) ;
    OBUF \out_obuf(394)  (.O (out[394]), .I (out_dup_0[394])) ;
    OBUF \out_obuf(395)  (.O (out[395]), .I (out_dup_0[395])) ;
    OBUF \out_obuf(396)  (.O (out[396]), .I (out_dup_0[396])) ;
    OBUF \out_obuf(397)  (.O (out[397]), .I (out_dup_0[397])) ;
    OBUF \out_obuf(398)  (.O (out[398]), .I (out_dup_0[398])) ;
    OBUF \out_obuf(399)  (.O (out[399]), .I (out_dup_0[399])) ;
    OBUF \out_obuf(400)  (.O (out[400]), .I (out_dup_0[400])) ;
    OBUF \out_obuf(401)  (.O (out[401]), .I (out_dup_0[401])) ;
    OBUF \out_obuf(402)  (.O (out[402]), .I (out_dup_0[402])) ;
    OBUF \out_obuf(403)  (.O (out[403]), .I (out_dup_0[403])) ;
    OBUF \out_obuf(404)  (.O (out[404]), .I (out_dup_0[404])) ;
    OBUF \out_obuf(405)  (.O (out[405]), .I (out_dup_0[405])) ;
    OBUF \out_obuf(406)  (.O (out[406]), .I (out_dup_0[406])) ;
    OBUF \out_obuf(407)  (.O (out[407]), .I (out_dup_0[407])) ;
    OBUF \out_obuf(408)  (.O (out[408]), .I (out_dup_0[408])) ;
    OBUF \out_obuf(409)  (.O (out[409]), .I (out_dup_0[409])) ;
    OBUF \out_obuf(410)  (.O (out[410]), .I (out_dup_0[410])) ;
    OBUF \out_obuf(411)  (.O (out[411]), .I (out_dup_0[411])) ;
    OBUF \out_obuf(412)  (.O (out[412]), .I (out_dup_0[412])) ;
    OBUF \out_obuf(413)  (.O (out[413]), .I (out_dup_0[413])) ;
    OBUF \out_obuf(414)  (.O (out[414]), .I (out_dup_0[414])) ;
    OBUF \out_obuf(415)  (.O (out[415]), .I (out_dup_0[415])) ;
    OBUF \out_obuf(416)  (.O (out[416]), .I (out_dup_0[416])) ;
    OBUF \out_obuf(417)  (.O (out[417]), .I (out_dup_0[417])) ;
    OBUF \out_obuf(418)  (.O (out[418]), .I (out_dup_0[418])) ;
    OBUF \out_obuf(419)  (.O (out[419]), .I (out_dup_0[419])) ;
    OBUF \out_obuf(420)  (.O (out[420]), .I (out_dup_0[420])) ;
    OBUF \out_obuf(421)  (.O (out[421]), .I (out_dup_0[421])) ;
    OBUF \out_obuf(422)  (.O (out[422]), .I (out_dup_0[422])) ;
    OBUF \out_obuf(423)  (.O (out[423]), .I (out_dup_0[423])) ;
    OBUF \out_obuf(424)  (.O (out[424]), .I (out_dup_0[424])) ;
    OBUF \out_obuf(425)  (.O (out[425]), .I (out_dup_0[425])) ;
    OBUF \out_obuf(426)  (.O (out[426]), .I (out_dup_0[426])) ;
    OBUF \out_obuf(427)  (.O (out[427]), .I (out_dup_0[427])) ;
    OBUF \out_obuf(428)  (.O (out[428]), .I (out_dup_0[428])) ;
    OBUF \out_obuf(429)  (.O (out[429]), .I (out_dup_0[429])) ;
    OBUF \out_obuf(430)  (.O (out[430]), .I (out_dup_0[430])) ;
    OBUF \out_obuf(431)  (.O (out[431]), .I (out_dup_0[431])) ;
    OBUF \out_obuf(432)  (.O (out[432]), .I (out_dup_0[432])) ;
    OBUF \out_obuf(433)  (.O (out[433]), .I (out_dup_0[433])) ;
    OBUF \out_obuf(434)  (.O (out[434]), .I (out_dup_0[434])) ;
    OBUF \out_obuf(435)  (.O (out[435]), .I (out_dup_0[435])) ;
    OBUF \out_obuf(436)  (.O (out[436]), .I (out_dup_0[436])) ;
    OBUF \out_obuf(437)  (.O (out[437]), .I (out_dup_0[437])) ;
    OBUF \out_obuf(438)  (.O (out[438]), .I (out_dup_0[438])) ;
    OBUF \out_obuf(439)  (.O (out[439]), .I (out_dup_0[439])) ;
    OBUF \out_obuf(440)  (.O (out[440]), .I (out_dup_0[440])) ;
    OBUF \out_obuf(441)  (.O (out[441]), .I (out_dup_0[441])) ;
    OBUF \out_obuf(442)  (.O (out[442]), .I (out_dup_0[442])) ;
    OBUF \out_obuf(443)  (.O (out[443]), .I (out_dup_0[443])) ;
    OBUF \out_obuf(444)  (.O (out[444]), .I (out_dup_0[444])) ;
    OBUF \out_obuf(445)  (.O (out[445]), .I (out_dup_0[445])) ;
    OBUF \out_obuf(446)  (.O (out[446]), .I (out_dup_0[446])) ;
    OBUF \out_obuf(447)  (.O (out[447]), .I (out_dup_0[447])) ;
    OBUF \out_obuf(448)  (.O (out[448]), .I (out_dup_0[448])) ;
    OBUF \out_obuf(449)  (.O (out[449]), .I (out_dup_0[449])) ;
    OBUF \out_obuf(450)  (.O (out[450]), .I (out_dup_0[450])) ;
    OBUF \out_obuf(451)  (.O (out[451]), .I (out_dup_0[451])) ;
    OBUF \out_obuf(452)  (.O (out[452]), .I (out_dup_0[452])) ;
    OBUF \out_obuf(453)  (.O (out[453]), .I (out_dup_0[453])) ;
    OBUF \out_obuf(454)  (.O (out[454]), .I (out_dup_0[454])) ;
    OBUF \out_obuf(455)  (.O (out[455]), .I (out_dup_0[455])) ;
    OBUF \out_obuf(456)  (.O (out[456]), .I (out_dup_0[456])) ;
    OBUF \out_obuf(457)  (.O (out[457]), .I (out_dup_0[457])) ;
    OBUF \out_obuf(458)  (.O (out[458]), .I (out_dup_0[458])) ;
    OBUF \out_obuf(459)  (.O (out[459]), .I (out_dup_0[459])) ;
    OBUF \out_obuf(460)  (.O (out[460]), .I (out_dup_0[460])) ;
    OBUF \out_obuf(461)  (.O (out[461]), .I (out_dup_0[461])) ;
    OBUF \out_obuf(462)  (.O (out[462]), .I (out_dup_0[462])) ;
    OBUF \out_obuf(463)  (.O (out[463]), .I (out_dup_0[463])) ;
    OBUF \out_obuf(464)  (.O (out[464]), .I (out_dup_0[464])) ;
    OBUF \out_obuf(465)  (.O (out[465]), .I (out_dup_0[465])) ;
    OBUF \out_obuf(466)  (.O (out[466]), .I (out_dup_0[466])) ;
    OBUF \out_obuf(467)  (.O (out[467]), .I (out_dup_0[467])) ;
    OBUF \out_obuf(468)  (.O (out[468]), .I (out_dup_0[468])) ;
    OBUF \out_obuf(469)  (.O (out[469]), .I (out_dup_0[469])) ;
    OBUF \out_obuf(470)  (.O (out[470]), .I (out_dup_0[470])) ;
    OBUF \out_obuf(471)  (.O (out[471]), .I (out_dup_0[471])) ;
    OBUF \out_obuf(472)  (.O (out[472]), .I (out_dup_0[472])) ;
    OBUF \out_obuf(473)  (.O (out[473]), .I (out_dup_0[473])) ;
    OBUF \out_obuf(474)  (.O (out[474]), .I (out_dup_0[474])) ;
    OBUF \out_obuf(475)  (.O (out[475]), .I (out_dup_0[475])) ;
    OBUF \out_obuf(476)  (.O (out[476]), .I (out_dup_0[476])) ;
    OBUF \out_obuf(477)  (.O (out[477]), .I (out_dup_0[477])) ;
    OBUF \out_obuf(478)  (.O (out[478]), .I (out_dup_0[478])) ;
    OBUF \out_obuf(479)  (.O (out[479]), .I (out_dup_0[479])) ;
    OBUF \out_obuf(480)  (.O (out[480]), .I (out_dup_0[480])) ;
    OBUF \out_obuf(481)  (.O (out[481]), .I (out_dup_0[481])) ;
    OBUF \out_obuf(482)  (.O (out[482]), .I (out_dup_0[482])) ;
    OBUF \out_obuf(483)  (.O (out[483]), .I (out_dup_0[483])) ;
    OBUF \out_obuf(484)  (.O (out[484]), .I (out_dup_0[484])) ;
    OBUF \out_obuf(485)  (.O (out[485]), .I (out_dup_0[485])) ;
    OBUF \out_obuf(486)  (.O (out[486]), .I (out_dup_0[486])) ;
    OBUF \out_obuf(487)  (.O (out[487]), .I (out_dup_0[487])) ;
    OBUF \out_obuf(488)  (.O (out[488]), .I (out_dup_0[488])) ;
    OBUF \out_obuf(489)  (.O (out[489]), .I (out_dup_0[489])) ;
    OBUF \out_obuf(490)  (.O (out[490]), .I (out_dup_0[490])) ;
    OBUF \out_obuf(491)  (.O (out[491]), .I (out_dup_0[491])) ;
    OBUF \out_obuf(492)  (.O (out[492]), .I (out_dup_0[492])) ;
    OBUF \out_obuf(493)  (.O (out[493]), .I (out_dup_0[493])) ;
    OBUF \out_obuf(494)  (.O (out[494]), .I (out_dup_0[494])) ;
    OBUF \out_obuf(495)  (.O (out[495]), .I (out_dup_0[495])) ;
    OBUF \out_obuf(496)  (.O (out[496]), .I (out_dup_0[496])) ;
    OBUF \out_obuf(497)  (.O (out[497]), .I (out_dup_0[497])) ;
    OBUF \out_obuf(498)  (.O (out[498]), .I (out_dup_0[498])) ;
    OBUF \out_obuf(499)  (.O (out[499]), .I (out_dup_0[499])) ;
    OBUF \out_obuf(500)  (.O (out[500]), .I (out_dup_0[500])) ;
    OBUF \out_obuf(501)  (.O (out[501]), .I (out_dup_0[501])) ;
    OBUF \out_obuf(502)  (.O (out[502]), .I (out_dup_0[502])) ;
    OBUF \out_obuf(503)  (.O (out[503]), .I (out_dup_0[503])) ;
    OBUF \out_obuf(504)  (.O (out[504]), .I (out_dup_0[504])) ;
    OBUF \out_obuf(505)  (.O (out[505]), .I (out_dup_0[505])) ;
    OBUF \out_obuf(506)  (.O (out[506]), .I (out_dup_0[506])) ;
    OBUF \out_obuf(507)  (.O (out[507]), .I (out_dup_0[507])) ;
    OBUF \out_obuf(508)  (.O (out[508]), .I (out_dup_0[508])) ;
    OBUF \out_obuf(509)  (.O (out[509]), .I (out_dup_0[509])) ;
    OBUF \out_obuf(510)  (.O (out[510]), .I (out_dup_0[510])) ;
    OBUF \out_obuf(511)  (.O (out[511]), .I (out_dup_0[511])) ;
    IBUF \in_ibuf(0)  (.O (in_int[70]), .I (in[0])) ;
    IBUF \in_ibuf(1)  (.O (in_int[71]), .I (in[1])) ;
    IBUF \in_ibuf(2)  (.O (in_int[72]), .I (in[2])) ;
    IBUF \in_ibuf(3)  (.O (in_int[73]), .I (in[3])) ;
    IBUF \in_ibuf(4)  (.O (in_int[74]), .I (in[4])) ;
    IBUF \in_ibuf(5)  (.O (in_int[75]), .I (in[5])) ;
    IBUF \in_ibuf(6)  (.O (in_int[76]), .I (in[6])) ;
    IBUF \in_ibuf(7)  (.O (in_int[77]), .I (in[7])) ;
    IBUF \in_ibuf(8)  (.O (in_int[78]), .I (in[8])) ;
    IBUF \in_ibuf(9)  (.O (in_int[79]), .I (in[9])) ;
    IBUF \in_ibuf(10)  (.O (in_int[80]), .I (in[10])) ;
    IBUF \in_ibuf(11)  (.O (in_int[81]), .I (in[11])) ;
    IBUF \in_ibuf(12)  (.O (in_int[82]), .I (in[12])) ;
    IBUF \in_ibuf(13)  (.O (in_int[83]), .I (in[13])) ;
    IBUF \in_ibuf(14)  (.O (in_int[84]), .I (in[14])) ;
    IBUF \in_ibuf(15)  (.O (in_int[85]), .I (in[15])) ;
    IBUF \in_ibuf(16)  (.O (in_int[86]), .I (in[16])) ;
    IBUF \in_ibuf(17)  (.O (in_int[87]), .I (in[17])) ;
    IBUF \in_ibuf(18)  (.O (in_int[88]), .I (in[18])) ;
    IBUF \in_ibuf(19)  (.O (in_int[89]), .I (in[19])) ;
    IBUF \in_ibuf(20)  (.O (in_int[90]), .I (in[20])) ;
    IBUF \in_ibuf(21)  (.O (in_int[91]), .I (in[21])) ;
    IBUF \in_ibuf(22)  (.O (in_int[92]), .I (in[22])) ;
    IBUF \in_ibuf(23)  (.O (in_int[93]), .I (in[23])) ;
    IBUF \in_ibuf(24)  (.O (in_int[94]), .I (in[24])) ;
    IBUF \in_ibuf(25)  (.O (in_int[95]), .I (in[25])) ;
    IBUF \in_ibuf(26)  (.O (in_int[96]), .I (in[26])) ;
    IBUF \in_ibuf(27)  (.O (in_int[97]), .I (in[27])) ;
    IBUF \in_ibuf(28)  (.O (in_int[98]), .I (in[28])) ;
    IBUF \in_ibuf(29)  (.O (in_int[99]), .I (in[29])) ;
    IBUF \in_ibuf(30)  (.O (in_int[100]), .I (in[30])) ;
    IBUF \in_ibuf(31)  (.O (in_int[101]), .I (in[31])) ;
    IBUF \in_ibuf(32)  (.O (in_int[102]), .I (in[32])) ;
    IBUF \in_ibuf(33)  (.O (in_int[103]), .I (in[33])) ;
    IBUF \in_ibuf(34)  (.O (in_int[104]), .I (in[34])) ;
    IBUF \in_ibuf(35)  (.O (in_int[105]), .I (in[35])) ;
    IBUF \in_ibuf(36)  (.O (in_int[106]), .I (in[36])) ;
    IBUF \in_ibuf(37)  (.O (in_int[107]), .I (in[37])) ;
    IBUF \in_ibuf(38)  (.O (in_int[108]), .I (in[38])) ;
    IBUF \in_ibuf(39)  (.O (in_int[109]), .I (in[39])) ;
    IBUF \in_ibuf(40)  (.O (in_int[110]), .I (in[40])) ;
    IBUF \in_ibuf(41)  (.O (in_int[111]), .I (in[41])) ;
    IBUF \in_ibuf(42)  (.O (in_int[112]), .I (in[42])) ;
    IBUF \in_ibuf(43)  (.O (in_int[113]), .I (in[43])) ;
    IBUF \in_ibuf(44)  (.O (in_int[114]), .I (in[44])) ;
    IBUF \in_ibuf(45)  (.O (in_int[115]), .I (in[45])) ;
    IBUF \in_ibuf(46)  (.O (in_int[116]), .I (in[46])) ;
    IBUF \in_ibuf(47)  (.O (in_int[117]), .I (in[47])) ;
    IBUF \in_ibuf(48)  (.O (in_int[118]), .I (in[48])) ;
    IBUF \in_ibuf(49)  (.O (in_int[119]), .I (in[49])) ;
    IBUF \in_ibuf(50)  (.O (in_int[120]), .I (in[50])) ;
    IBUF \in_ibuf(51)  (.O (in_int[121]), .I (in[51])) ;
    IBUF \in_ibuf(52)  (.O (in_int[122]), .I (in[52])) ;
    IBUF \in_ibuf(53)  (.O (in_int[123]), .I (in[53])) ;
    IBUF \in_ibuf(54)  (.O (in_int[124]), .I (in[54])) ;
    IBUF \in_ibuf(55)  (.O (in_int[125]), .I (in[55])) ;
    IBUF \in_ibuf(56)  (.O (in_int[126]), .I (in[56])) ;
    IBUF \in_ibuf(57)  (.O (in_int[127]), .I (in[57])) ;
    IBUF \in_ibuf(58)  (.O (in_int[128]), .I (in[58])) ;
    IBUF \in_ibuf(59)  (.O (in_int[129]), .I (in[59])) ;
    IBUF \in_ibuf(60)  (.O (in_int[130]), .I (in[60])) ;
    IBUF \in_ibuf(61)  (.O (in_int[131]), .I (in[61])) ;
    IBUF \in_ibuf(62)  (.O (in_int[132]), .I (in[62])) ;
    IBUF \in_ibuf(63)  (.O (in_int[133]), .I (in[63])) ;
    IBUF \in_ibuf(64)  (.O (in_int[134]), .I (in[64])) ;
    IBUF \in_ibuf(65)  (.O (in_int[135]), .I (in[65])) ;
    IBUF \in_ibuf(66)  (.O (in_int[136]), .I (in[66])) ;
    IBUF \in_ibuf(67)  (.O (in_int[137]), .I (in[67])) ;
    IBUF \in_ibuf(68)  (.O (in_int[138]), .I (in[68])) ;
    IBUF \in_ibuf(69)  (.O (in_int[139]), .I (in[69])) ;
    IBUF \in_ibuf(70)  (.O (in_int[140]), .I (in[70])) ;
    IBUF \in_ibuf(71)  (.O (in_int[141]), .I (in[71])) ;
    IBUF \in_ibuf(72)  (.O (in_int[142]), .I (in[72])) ;
    IBUF \in_ibuf(73)  (.O (in_int[143]), .I (in[73])) ;
    IBUF \in_ibuf(74)  (.O (in_int[144]), .I (in[74])) ;
    IBUF \in_ibuf(75)  (.O (in_int[145]), .I (in[75])) ;
    IBUF \in_ibuf(76)  (.O (in_int[146]), .I (in[76])) ;
    IBUF \in_ibuf(77)  (.O (in_int[147]), .I (in[77])) ;
    IBUF \in_ibuf(78)  (.O (in_int[148]), .I (in[78])) ;
    IBUF \in_ibuf(79)  (.O (in_int[149]), .I (in[79])) ;
    IBUF \in_ibuf(80)  (.O (in_int[150]), .I (in[80])) ;
    IBUF \in_ibuf(81)  (.O (in_int[151]), .I (in[81])) ;
    IBUF \in_ibuf(82)  (.O (in_int[152]), .I (in[82])) ;
    IBUF \in_ibuf(83)  (.O (in_int[153]), .I (in[83])) ;
    IBUF \in_ibuf(84)  (.O (in_int[154]), .I (in[84])) ;
    IBUF \in_ibuf(85)  (.O (in_int[155]), .I (in[85])) ;
    IBUF \in_ibuf(86)  (.O (in_int[156]), .I (in[86])) ;
    IBUF \in_ibuf(87)  (.O (in_int[157]), .I (in[87])) ;
    IBUF \in_ibuf(88)  (.O (in_int[158]), .I (in[88])) ;
    IBUF \in_ibuf(89)  (.O (in_int[159]), .I (in[89])) ;
    IBUF \in_ibuf(90)  (.O (in_int[160]), .I (in[90])) ;
    IBUF \in_ibuf(91)  (.O (in_int[161]), .I (in[91])) ;
    IBUF \in_ibuf(92)  (.O (in_int[162]), .I (in[92])) ;
    IBUF \in_ibuf(93)  (.O (in_int[163]), .I (in[93])) ;
    IBUF \in_ibuf(94)  (.O (in_int[164]), .I (in[94])) ;
    IBUF \in_ibuf(95)  (.O (in_int[165]), .I (in[95])) ;
    IBUF \in_ibuf(96)  (.O (in_int[166]), .I (in[96])) ;
    IBUF \in_ibuf(97)  (.O (in_int[167]), .I (in[97])) ;
    IBUF \in_ibuf(98)  (.O (in_int[168]), .I (in[98])) ;
    IBUF \in_ibuf(99)  (.O (in_int[169]), .I (in[99])) ;
    IBUF \in_ibuf(100)  (.O (in_int[170]), .I (in[100])) ;
    IBUF \in_ibuf(101)  (.O (in_int[171]), .I (in[101])) ;
    IBUF \in_ibuf(102)  (.O (in_int[172]), .I (in[102])) ;
    IBUF \in_ibuf(103)  (.O (in_int[173]), .I (in[103])) ;
    IBUF \in_ibuf(104)  (.O (in_int[174]), .I (in[104])) ;
    IBUF \in_ibuf(105)  (.O (in_int[175]), .I (in[105])) ;
    IBUF \in_ibuf(106)  (.O (in_int[176]), .I (in[106])) ;
    IBUF \in_ibuf(107)  (.O (in_int[177]), .I (in[107])) ;
    IBUF \in_ibuf(108)  (.O (in_int[178]), .I (in[108])) ;
    IBUF \in_ibuf(109)  (.O (in_int[179]), .I (in[109])) ;
    IBUF \in_ibuf(110)  (.O (in_int[180]), .I (in[110])) ;
    IBUF \in_ibuf(111)  (.O (in_int[181]), .I (in[111])) ;
    IBUF \in_ibuf(112)  (.O (in_int[182]), .I (in[112])) ;
    IBUF \in_ibuf(113)  (.O (in_int[183]), .I (in[113])) ;
    IBUF \in_ibuf(114)  (.O (in_int[184]), .I (in[114])) ;
    IBUF \in_ibuf(115)  (.O (in_int[185]), .I (in[115])) ;
    IBUF \in_ibuf(116)  (.O (in_int[186]), .I (in[116])) ;
    IBUF \in_ibuf(117)  (.O (in_int[187]), .I (in[117])) ;
    IBUF \in_ibuf(118)  (.O (in_int[188]), .I (in[118])) ;
    IBUF \in_ibuf(119)  (.O (in_int[189]), .I (in[119])) ;
    IBUF \in_ibuf(120)  (.O (in_int[190]), .I (in[120])) ;
    IBUF \in_ibuf(121)  (.O (in_int[191]), .I (in[121])) ;
    IBUF \in_ibuf(122)  (.O (in_int[192]), .I (in[122])) ;
    IBUF \in_ibuf(123)  (.O (in_int[193]), .I (in[123])) ;
    IBUF \in_ibuf(124)  (.O (in_int[194]), .I (in[124])) ;
    IBUF \in_ibuf(125)  (.O (in_int[195]), .I (in[125])) ;
    IBUF \in_ibuf(126)  (.O (in_int[196]), .I (in[126])) ;
    IBUF \in_ibuf(127)  (.O (in_int[197]), .I (in[127])) ;
    IBUF \in_ibuf(128)  (.O (in_int[198]), .I (in[128])) ;
    IBUF \in_ibuf(129)  (.O (in_int[199]), .I (in[129])) ;
    IBUF \in_ibuf(130)  (.O (in_int[200]), .I (in[130])) ;
    IBUF \in_ibuf(131)  (.O (in_int[201]), .I (in[131])) ;
    IBUF \in_ibuf(132)  (.O (in_int[202]), .I (in[132])) ;
    IBUF \in_ibuf(133)  (.O (in_int[203]), .I (in[133])) ;
    IBUF \in_ibuf(134)  (.O (in_int[204]), .I (in[134])) ;
    IBUF \in_ibuf(135)  (.O (in_int[205]), .I (in[135])) ;
    IBUF \in_ibuf(136)  (.O (in_int[206]), .I (in[136])) ;
    IBUF \in_ibuf(137)  (.O (in_int[207]), .I (in[137])) ;
    IBUF \in_ibuf(138)  (.O (in_int[208]), .I (in[138])) ;
    IBUF \in_ibuf(139)  (.O (in_int[209]), .I (in[139])) ;
    IBUF \in_ibuf(140)  (.O (in_int[210]), .I (in[140])) ;
    IBUF \in_ibuf(141)  (.O (in_int[211]), .I (in[141])) ;
    IBUF \in_ibuf(142)  (.O (in_int[212]), .I (in[142])) ;
    IBUF \in_ibuf(143)  (.O (in_int[213]), .I (in[143])) ;
    IBUF \in_ibuf(144)  (.O (in_int[214]), .I (in[144])) ;
    IBUF \in_ibuf(145)  (.O (in_int[215]), .I (in[145])) ;
    IBUF \in_ibuf(146)  (.O (in_int[216]), .I (in[146])) ;
    IBUF \in_ibuf(147)  (.O (in_int[217]), .I (in[147])) ;
    IBUF \in_ibuf(148)  (.O (in_int[218]), .I (in[148])) ;
    IBUF \in_ibuf(149)  (.O (in_int[219]), .I (in[149])) ;
    IBUF \in_ibuf(150)  (.O (in_int[220]), .I (in[150])) ;
    IBUF \in_ibuf(151)  (.O (in_int[221]), .I (in[151])) ;
    IBUF \in_ibuf(152)  (.O (in_int[222]), .I (in[152])) ;
    IBUF \in_ibuf(153)  (.O (in_int[223]), .I (in[153])) ;
    IBUF \in_ibuf(154)  (.O (in_int[224]), .I (in[154])) ;
    IBUF \in_ibuf(155)  (.O (in_int[225]), .I (in[155])) ;
    IBUF \in_ibuf(156)  (.O (in_int[226]), .I (in[156])) ;
    IBUF \in_ibuf(157)  (.O (in_int[227]), .I (in[157])) ;
    IBUF \in_ibuf(158)  (.O (in_int[228]), .I (in[158])) ;
    IBUF \in_ibuf(159)  (.O (in_int[229]), .I (in[159])) ;
    IBUF \in_ibuf(160)  (.O (in_int[230]), .I (in[160])) ;
    IBUF \in_ibuf(161)  (.O (in_int[231]), .I (in[161])) ;
    IBUF \in_ibuf(162)  (.O (in_int[232]), .I (in[162])) ;
    IBUF \in_ibuf(163)  (.O (in_int[233]), .I (in[163])) ;
    IBUF \in_ibuf(164)  (.O (in_int[234]), .I (in[164])) ;
    IBUF \in_ibuf(165)  (.O (in_int[235]), .I (in[165])) ;
    IBUF \in_ibuf(166)  (.O (in_int[236]), .I (in[166])) ;
    IBUF \in_ibuf(167)  (.O (in_int[237]), .I (in[167])) ;
    IBUF \in_ibuf(168)  (.O (in_int[238]), .I (in[168])) ;
    IBUF \in_ibuf(169)  (.O (in_int[239]), .I (in[169])) ;
    IBUF \in_ibuf(170)  (.O (in_int[240]), .I (in[170])) ;
    IBUF \in_ibuf(171)  (.O (in_int[241]), .I (in[171])) ;
    IBUF \in_ibuf(172)  (.O (in_int[242]), .I (in[172])) ;
    IBUF \in_ibuf(173)  (.O (in_int[243]), .I (in[173])) ;
    IBUF \in_ibuf(174)  (.O (in_int[244]), .I (in[174])) ;
    IBUF \in_ibuf(175)  (.O (in_int[245]), .I (in[175])) ;
    IBUF \in_ibuf(176)  (.O (in_int[246]), .I (in[176])) ;
    IBUF \in_ibuf(177)  (.O (in_int[247]), .I (in[177])) ;
    IBUF \in_ibuf(178)  (.O (in_int[248]), .I (in[178])) ;
    IBUF \in_ibuf(179)  (.O (in_int[249]), .I (in[179])) ;
    IBUF \in_ibuf(180)  (.O (in_int[250]), .I (in[180])) ;
    IBUF \in_ibuf(181)  (.O (in_int[251]), .I (in[181])) ;
    IBUF \in_ibuf(182)  (.O (in_int[252]), .I (in[182])) ;
    IBUF \in_ibuf(183)  (.O (in_int[253]), .I (in[183])) ;
    IBUF \in_ibuf(184)  (.O (in_int[254]), .I (in[184])) ;
    IBUF \in_ibuf(185)  (.O (in_int[255]), .I (in[185])) ;
    IBUF \in_ibuf(186)  (.O (in_int[256]), .I (in[186])) ;
    IBUF \in_ibuf(187)  (.O (in_int[257]), .I (in[187])) ;
    IBUF \in_ibuf(188)  (.O (in_int[258]), .I (in[188])) ;
    IBUF \in_ibuf(189)  (.O (in_int[259]), .I (in[189])) ;
    IBUF \in_ibuf(190)  (.O (in_int[260]), .I (in[190])) ;
    IBUF \in_ibuf(191)  (.O (in_int[261]), .I (in[191])) ;
    IBUF \in_ibuf(192)  (.O (in_int[262]), .I (in[192])) ;
    IBUF \in_ibuf(193)  (.O (in_int[263]), .I (in[193])) ;
    IBUF \in_ibuf(194)  (.O (in_int[264]), .I (in[194])) ;
    IBUF \in_ibuf(195)  (.O (in_int[265]), .I (in[195])) ;
    IBUF \in_ibuf(196)  (.O (in_int[266]), .I (in[196])) ;
    IBUF \in_ibuf(197)  (.O (in_int[267]), .I (in[197])) ;
    IBUF \in_ibuf(198)  (.O (in_int[268]), .I (in[198])) ;
    IBUF \in_ibuf(199)  (.O (in_int[269]), .I (in[199])) ;
    IBUF \in_ibuf(200)  (.O (in_int[270]), .I (in[200])) ;
    IBUF \in_ibuf(201)  (.O (in_int[271]), .I (in[201])) ;
    IBUF \in_ibuf(202)  (.O (in_int[272]), .I (in[202])) ;
    IBUF \in_ibuf(203)  (.O (in_int[273]), .I (in[203])) ;
    IBUF \in_ibuf(204)  (.O (in_int[274]), .I (in[204])) ;
    IBUF \in_ibuf(205)  (.O (in_int[275]), .I (in[205])) ;
    IBUF \in_ibuf(206)  (.O (in_int[276]), .I (in[206])) ;
    IBUF \in_ibuf(207)  (.O (in_int[277]), .I (in[207])) ;
    IBUF \in_ibuf(208)  (.O (in_int[278]), .I (in[208])) ;
    IBUF \in_ibuf(209)  (.O (in_int[279]), .I (in[209])) ;
    IBUF \in_ibuf(210)  (.O (in_int[280]), .I (in[210])) ;
    IBUF \in_ibuf(211)  (.O (in_int[281]), .I (in[211])) ;
    IBUF \in_ibuf(212)  (.O (in_int[282]), .I (in[212])) ;
    IBUF \in_ibuf(213)  (.O (in_int[283]), .I (in[213])) ;
    IBUF \in_ibuf(214)  (.O (in_int[284]), .I (in[214])) ;
    IBUF \in_ibuf(215)  (.O (in_int[285]), .I (in[215])) ;
    IBUF \in_ibuf(216)  (.O (in_int[286]), .I (in[216])) ;
    IBUF \in_ibuf(217)  (.O (in_int[287]), .I (in[217])) ;
    IBUF \in_ibuf(218)  (.O (in_int[288]), .I (in[218])) ;
    IBUF \in_ibuf(219)  (.O (in_int[289]), .I (in[219])) ;
    IBUF \in_ibuf(220)  (.O (in_int[290]), .I (in[220])) ;
    IBUF \in_ibuf(221)  (.O (in_int[291]), .I (in[221])) ;
    IBUF \in_ibuf(222)  (.O (in_int[292]), .I (in[222])) ;
    IBUF \in_ibuf(223)  (.O (in_int[293]), .I (in[223])) ;
    IBUF \in_ibuf(224)  (.O (in_int[294]), .I (in[224])) ;
    IBUF \in_ibuf(225)  (.O (in_int[295]), .I (in[225])) ;
    IBUF \in_ibuf(226)  (.O (in_int[296]), .I (in[226])) ;
    IBUF \in_ibuf(227)  (.O (in_int[297]), .I (in[227])) ;
    IBUF \in_ibuf(228)  (.O (in_int[298]), .I (in[228])) ;
    IBUF \in_ibuf(229)  (.O (in_int[299]), .I (in[229])) ;
    IBUF \in_ibuf(230)  (.O (in_int[300]), .I (in[230])) ;
    IBUF \in_ibuf(231)  (.O (in_int[301]), .I (in[231])) ;
    IBUF \in_ibuf(232)  (.O (in_int[302]), .I (in[232])) ;
    IBUF \in_ibuf(233)  (.O (in_int[303]), .I (in[233])) ;
    IBUF \in_ibuf(234)  (.O (in_int[304]), .I (in[234])) ;
    IBUF \in_ibuf(235)  (.O (in_int[305]), .I (in[235])) ;
    IBUF \in_ibuf(236)  (.O (in_int[306]), .I (in[236])) ;
    IBUF \in_ibuf(237)  (.O (in_int[307]), .I (in[237])) ;
    IBUF \in_ibuf(238)  (.O (in_int[308]), .I (in[238])) ;
    IBUF \in_ibuf(239)  (.O (in_int[309]), .I (in[239])) ;
    IBUF \in_ibuf(240)  (.O (in_int[310]), .I (in[240])) ;
    IBUF \in_ibuf(241)  (.O (in_int[311]), .I (in[241])) ;
    IBUF \in_ibuf(242)  (.O (in_int[312]), .I (in[242])) ;
    IBUF \in_ibuf(243)  (.O (in_int[313]), .I (in[243])) ;
    IBUF \in_ibuf(244)  (.O (in_int[314]), .I (in[244])) ;
    IBUF \in_ibuf(245)  (.O (in_int[315]), .I (in[245])) ;
    IBUF \in_ibuf(246)  (.O (in_int[316]), .I (in[246])) ;
    IBUF \in_ibuf(247)  (.O (in_int[317]), .I (in[247])) ;
    IBUF \in_ibuf(248)  (.O (in_int[318]), .I (in[248])) ;
    IBUF \in_ibuf(249)  (.O (in_int[319]), .I (in[249])) ;
    IBUF \in_ibuf(250)  (.O (in_int[320]), .I (in[250])) ;
    IBUF \in_ibuf(251)  (.O (in_int[321]), .I (in[251])) ;
    IBUF \in_ibuf(252)  (.O (in_int[322]), .I (in[252])) ;
    IBUF \in_ibuf(253)  (.O (in_int[323]), .I (in[253])) ;
    IBUF \in_ibuf(254)  (.O (in_int[324]), .I (in[254])) ;
    IBUF \in_ibuf(255)  (.O (in_int[325]), .I (in[255])) ;
    IBUF \in_ibuf(256)  (.O (in_int[326]), .I (in[256])) ;
    IBUF \in_ibuf(257)  (.O (in_int[327]), .I (in[257])) ;
    IBUF \in_ibuf(258)  (.O (in_int[328]), .I (in[258])) ;
    IBUF \in_ibuf(259)  (.O (in_int[329]), .I (in[259])) ;
    IBUF \in_ibuf(260)  (.O (in_int[330]), .I (in[260])) ;
    IBUF \in_ibuf(261)  (.O (in_int[331]), .I (in[261])) ;
    IBUF \in_ibuf(262)  (.O (in_int[332]), .I (in[262])) ;
    IBUF \in_ibuf(263)  (.O (in_int[333]), .I (in[263])) ;
    IBUF \in_ibuf(264)  (.O (in_int[334]), .I (in[264])) ;
    IBUF \in_ibuf(265)  (.O (in_int[335]), .I (in[265])) ;
    IBUF \in_ibuf(266)  (.O (in_int[336]), .I (in[266])) ;
    IBUF \in_ibuf(267)  (.O (in_int[337]), .I (in[267])) ;
    IBUF \in_ibuf(268)  (.O (in_int[338]), .I (in[268])) ;
    IBUF \in_ibuf(269)  (.O (in_int[339]), .I (in[269])) ;
    IBUF \in_ibuf(270)  (.O (in_int[340]), .I (in[270])) ;
    IBUF \in_ibuf(271)  (.O (in_int[341]), .I (in[271])) ;
    IBUF \in_ibuf(272)  (.O (in_int[342]), .I (in[272])) ;
    IBUF \in_ibuf(273)  (.O (in_int[343]), .I (in[273])) ;
    IBUF \in_ibuf(274)  (.O (in_int[344]), .I (in[274])) ;
    IBUF \in_ibuf(275)  (.O (in_int[345]), .I (in[275])) ;
    IBUF \in_ibuf(276)  (.O (in_int[346]), .I (in[276])) ;
    IBUF \in_ibuf(277)  (.O (in_int[347]), .I (in[277])) ;
    IBUF \in_ibuf(278)  (.O (in_int[348]), .I (in[278])) ;
    IBUF \in_ibuf(279)  (.O (in_int[349]), .I (in[279])) ;
    IBUF \in_ibuf(280)  (.O (in_int[350]), .I (in[280])) ;
    IBUF \in_ibuf(281)  (.O (in_int[351]), .I (in[281])) ;
    IBUF \in_ibuf(282)  (.O (in_int[352]), .I (in[282])) ;
    IBUF \in_ibuf(283)  (.O (in_int[353]), .I (in[283])) ;
    IBUF \in_ibuf(284)  (.O (in_int[354]), .I (in[284])) ;
    IBUF \in_ibuf(285)  (.O (in_int[355]), .I (in[285])) ;
    IBUF \in_ibuf(286)  (.O (in_int[356]), .I (in[286])) ;
    IBUF \in_ibuf(287)  (.O (in_int[357]), .I (in[287])) ;
    IBUF \in_ibuf(288)  (.O (in_int[358]), .I (in[288])) ;
    IBUF \in_ibuf(289)  (.O (in_int[359]), .I (in[289])) ;
    IBUF \in_ibuf(290)  (.O (in_int[360]), .I (in[290])) ;
    IBUF \in_ibuf(291)  (.O (in_int[361]), .I (in[291])) ;
    IBUF \in_ibuf(292)  (.O (in_int[362]), .I (in[292])) ;
    IBUF \in_ibuf(293)  (.O (in_int[363]), .I (in[293])) ;
    IBUF \in_ibuf(294)  (.O (in_int[364]), .I (in[294])) ;
    IBUF \in_ibuf(295)  (.O (in_int[365]), .I (in[295])) ;
    IBUF \in_ibuf(296)  (.O (in_int[366]), .I (in[296])) ;
    IBUF \in_ibuf(297)  (.O (in_int[367]), .I (in[297])) ;
    IBUF \in_ibuf(298)  (.O (in_int[368]), .I (in[298])) ;
    IBUF \in_ibuf(299)  (.O (in_int[369]), .I (in[299])) ;
    IBUF \in_ibuf(300)  (.O (in_int[370]), .I (in[300])) ;
    IBUF \in_ibuf(301)  (.O (in_int[371]), .I (in[301])) ;
    IBUF \in_ibuf(302)  (.O (in_int[372]), .I (in[302])) ;
    IBUF \in_ibuf(303)  (.O (in_int[373]), .I (in[303])) ;
    IBUF \in_ibuf(304)  (.O (in_int[374]), .I (in[304])) ;
    IBUF \in_ibuf(305)  (.O (in_int[375]), .I (in[305])) ;
    IBUF \in_ibuf(306)  (.O (in_int[376]), .I (in[306])) ;
    IBUF \in_ibuf(307)  (.O (in_int[377]), .I (in[307])) ;
    IBUF \in_ibuf(308)  (.O (in_int[378]), .I (in[308])) ;
    IBUF \in_ibuf(309)  (.O (in_int[379]), .I (in[309])) ;
    IBUF \in_ibuf(310)  (.O (in_int[380]), .I (in[310])) ;
    IBUF \in_ibuf(311)  (.O (in_int[381]), .I (in[311])) ;
    IBUF \in_ibuf(312)  (.O (in_int[382]), .I (in[312])) ;
    IBUF \in_ibuf(313)  (.O (in_int[383]), .I (in[313])) ;
    IBUF \in_ibuf(314)  (.O (in_int[384]), .I (in[314])) ;
    IBUF \in_ibuf(315)  (.O (in_int[385]), .I (in[315])) ;
    IBUF \in_ibuf(316)  (.O (in_int[386]), .I (in[316])) ;
    IBUF \in_ibuf(317)  (.O (in_int[387]), .I (in[317])) ;
    IBUF \in_ibuf(318)  (.O (in_int[388]), .I (in[318])) ;
    IBUF \in_ibuf(319)  (.O (in_int[389]), .I (in[319])) ;
    IBUF \in_ibuf(320)  (.O (in_int[390]), .I (in[320])) ;
    IBUF \in_ibuf(321)  (.O (in_int[391]), .I (in[321])) ;
    IBUF \in_ibuf(322)  (.O (in_int[392]), .I (in[322])) ;
    IBUF \in_ibuf(323)  (.O (in_int[393]), .I (in[323])) ;
    IBUF \in_ibuf(324)  (.O (in_int[394]), .I (in[324])) ;
    IBUF \in_ibuf(325)  (.O (in_int[395]), .I (in[325])) ;
    IBUF \in_ibuf(326)  (.O (in_int[396]), .I (in[326])) ;
    IBUF \in_ibuf(327)  (.O (in_int[397]), .I (in[327])) ;
    IBUF \in_ibuf(328)  (.O (in_int[398]), .I (in[328])) ;
    IBUF \in_ibuf(329)  (.O (in_int[399]), .I (in[329])) ;
    IBUF \in_ibuf(330)  (.O (in_int[400]), .I (in[330])) ;
    IBUF \in_ibuf(331)  (.O (in_int[401]), .I (in[331])) ;
    IBUF \in_ibuf(332)  (.O (in_int[402]), .I (in[332])) ;
    IBUF \in_ibuf(333)  (.O (in_int[403]), .I (in[333])) ;
    IBUF \in_ibuf(334)  (.O (in_int[404]), .I (in[334])) ;
    IBUF \in_ibuf(335)  (.O (in_int[405]), .I (in[335])) ;
    IBUF \in_ibuf(336)  (.O (in_int[406]), .I (in[336])) ;
    IBUF \in_ibuf(337)  (.O (in_int[407]), .I (in[337])) ;
    IBUF \in_ibuf(338)  (.O (in_int[408]), .I (in[338])) ;
    IBUF \in_ibuf(339)  (.O (in_int[409]), .I (in[339])) ;
    IBUF \in_ibuf(340)  (.O (in_int[410]), .I (in[340])) ;
    IBUF \in_ibuf(341)  (.O (in_int[411]), .I (in[341])) ;
    IBUF \in_ibuf(342)  (.O (in_int[412]), .I (in[342])) ;
    IBUF \in_ibuf(343)  (.O (in_int[413]), .I (in[343])) ;
    IBUF \in_ibuf(344)  (.O (in_int[414]), .I (in[344])) ;
    IBUF \in_ibuf(345)  (.O (in_int[415]), .I (in[345])) ;
    IBUF \in_ibuf(346)  (.O (in_int[416]), .I (in[346])) ;
    IBUF \in_ibuf(347)  (.O (in_int[417]), .I (in[347])) ;
    IBUF \in_ibuf(348)  (.O (in_int[418]), .I (in[348])) ;
    IBUF \in_ibuf(349)  (.O (in_int[419]), .I (in[349])) ;
    IBUF \in_ibuf(350)  (.O (in_int[420]), .I (in[350])) ;
    IBUF \in_ibuf(351)  (.O (in_int[421]), .I (in[351])) ;
    IBUF \in_ibuf(352)  (.O (in_int[422]), .I (in[352])) ;
    IBUF \in_ibuf(353)  (.O (in_int[423]), .I (in[353])) ;
    IBUF \in_ibuf(354)  (.O (in_int[424]), .I (in[354])) ;
    IBUF \in_ibuf(355)  (.O (in_int[425]), .I (in[355])) ;
    IBUF \in_ibuf(356)  (.O (in_int[426]), .I (in[356])) ;
    IBUF \in_ibuf(357)  (.O (in_int[427]), .I (in[357])) ;
    IBUF \in_ibuf(358)  (.O (in_int[428]), .I (in[358])) ;
    IBUF \in_ibuf(359)  (.O (in_int[429]), .I (in[359])) ;
    IBUF \in_ibuf(360)  (.O (in_int[430]), .I (in[360])) ;
    IBUF \in_ibuf(361)  (.O (in_int[431]), .I (in[361])) ;
    IBUF \in_ibuf(362)  (.O (in_int[432]), .I (in[362])) ;
    IBUF \in_ibuf(363)  (.O (in_int[433]), .I (in[363])) ;
    IBUF \in_ibuf(364)  (.O (in_int[434]), .I (in[364])) ;
    IBUF \in_ibuf(365)  (.O (in_int[435]), .I (in[365])) ;
    IBUF \in_ibuf(366)  (.O (in_int[436]), .I (in[366])) ;
    IBUF \in_ibuf(367)  (.O (in_int[437]), .I (in[367])) ;
    IBUF \in_ibuf(368)  (.O (in_int[438]), .I (in[368])) ;
    IBUF \in_ibuf(369)  (.O (in_int[439]), .I (in[369])) ;
    IBUF \in_ibuf(370)  (.O (in_int[440]), .I (in[370])) ;
    IBUF \in_ibuf(371)  (.O (in_int[441]), .I (in[371])) ;
    IBUF \in_ibuf(372)  (.O (in_int[442]), .I (in[372])) ;
    IBUF \in_ibuf(373)  (.O (in_int[443]), .I (in[373])) ;
    IBUF \in_ibuf(374)  (.O (in_int[444]), .I (in[374])) ;
    IBUF \in_ibuf(375)  (.O (in_int[445]), .I (in[375])) ;
    IBUF \in_ibuf(376)  (.O (in_int[446]), .I (in[376])) ;
    IBUF \in_ibuf(377)  (.O (in_int[447]), .I (in[377])) ;
    IBUF \in_ibuf(378)  (.O (in_int[448]), .I (in[378])) ;
    IBUF \in_ibuf(379)  (.O (in_int[449]), .I (in[379])) ;
    IBUF \in_ibuf(380)  (.O (in_int[450]), .I (in[380])) ;
    IBUF \in_ibuf(381)  (.O (in_int[451]), .I (in[381])) ;
    IBUF \in_ibuf(382)  (.O (in_int[452]), .I (in[382])) ;
    IBUF \in_ibuf(383)  (.O (in_int[453]), .I (in[383])) ;
    IBUF \in_ibuf(384)  (.O (in_int[454]), .I (in[384])) ;
    IBUF \in_ibuf(385)  (.O (in_int[455]), .I (in[385])) ;
    IBUF \in_ibuf(386)  (.O (in_int[456]), .I (in[386])) ;
    IBUF \in_ibuf(387)  (.O (in_int[457]), .I (in[387])) ;
    IBUF \in_ibuf(388)  (.O (in_int[458]), .I (in[388])) ;
    IBUF \in_ibuf(389)  (.O (in_int[459]), .I (in[389])) ;
    IBUF \in_ibuf(390)  (.O (in_int[460]), .I (in[390])) ;
    IBUF \in_ibuf(391)  (.O (in_int[461]), .I (in[391])) ;
    IBUF \in_ibuf(392)  (.O (in_int[462]), .I (in[392])) ;
    IBUF \in_ibuf(393)  (.O (in_int[463]), .I (in[393])) ;
    IBUF \in_ibuf(394)  (.O (in_int[464]), .I (in[394])) ;
    IBUF \in_ibuf(395)  (.O (in_int[465]), .I (in[395])) ;
    IBUF \in_ibuf(396)  (.O (in_int[466]), .I (in[396])) ;
    IBUF \in_ibuf(397)  (.O (in_int[467]), .I (in[397])) ;
    IBUF \in_ibuf(398)  (.O (in_int[468]), .I (in[398])) ;
    IBUF \in_ibuf(399)  (.O (in_int[469]), .I (in[399])) ;
    IBUF \in_ibuf(400)  (.O (in_int[470]), .I (in[400])) ;
    IBUF \in_ibuf(401)  (.O (in_int[471]), .I (in[401])) ;
    IBUF \in_ibuf(402)  (.O (in_int[472]), .I (in[402])) ;
    IBUF \in_ibuf(403)  (.O (in_int[473]), .I (in[403])) ;
    IBUF \in_ibuf(404)  (.O (in_int[474]), .I (in[404])) ;
    IBUF \in_ibuf(405)  (.O (in_int[475]), .I (in[405])) ;
    IBUF \in_ibuf(406)  (.O (in_int[476]), .I (in[406])) ;
    IBUF \in_ibuf(407)  (.O (in_int[477]), .I (in[407])) ;
    IBUF \in_ibuf(408)  (.O (in_int[478]), .I (in[408])) ;
    IBUF \in_ibuf(409)  (.O (in_int[479]), .I (in[409])) ;
    IBUF \in_ibuf(410)  (.O (in_int[480]), .I (in[410])) ;
    IBUF \in_ibuf(411)  (.O (in_int[481]), .I (in[411])) ;
    IBUF \in_ibuf(412)  (.O (in_int[482]), .I (in[412])) ;
    IBUF \in_ibuf(413)  (.O (in_int[483]), .I (in[413])) ;
    IBUF \in_ibuf(414)  (.O (in_int[484]), .I (in[414])) ;
    IBUF \in_ibuf(415)  (.O (in_int[485]), .I (in[415])) ;
    IBUF \in_ibuf(416)  (.O (in_int[486]), .I (in[416])) ;
    IBUF \in_ibuf(417)  (.O (in_int[487]), .I (in[417])) ;
    IBUF \in_ibuf(418)  (.O (in_int[488]), .I (in[418])) ;
    IBUF \in_ibuf(419)  (.O (in_int[489]), .I (in[419])) ;
    IBUF \in_ibuf(420)  (.O (in_int[490]), .I (in[420])) ;
    IBUF \in_ibuf(421)  (.O (in_int[491]), .I (in[421])) ;
    IBUF \in_ibuf(422)  (.O (in_int[492]), .I (in[422])) ;
    IBUF \in_ibuf(423)  (.O (in_int[493]), .I (in[423])) ;
    IBUF \in_ibuf(424)  (.O (in_int[494]), .I (in[424])) ;
    IBUF \in_ibuf(425)  (.O (in_int[495]), .I (in[425])) ;
    IBUF \in_ibuf(426)  (.O (in_int[496]), .I (in[426])) ;
    IBUF \in_ibuf(427)  (.O (in_int[497]), .I (in[427])) ;
    IBUF \in_ibuf(428)  (.O (in_int[498]), .I (in[428])) ;
    IBUF \in_ibuf(429)  (.O (in_int[499]), .I (in[429])) ;
    IBUF \in_ibuf(430)  (.O (in_int[500]), .I (in[430])) ;
    IBUF \in_ibuf(431)  (.O (in_int[501]), .I (in[431])) ;
    IBUF \in_ibuf(432)  (.O (in_int[502]), .I (in[432])) ;
    IBUF \in_ibuf(433)  (.O (in_int[503]), .I (in[433])) ;
    IBUF \in_ibuf(434)  (.O (in_int[504]), .I (in[434])) ;
    IBUF \in_ibuf(435)  (.O (in_int[505]), .I (in[435])) ;
    IBUF \in_ibuf(436)  (.O (in_int[506]), .I (in[436])) ;
    IBUF \in_ibuf(437)  (.O (in_int[507]), .I (in[437])) ;
    IBUF \in_ibuf(438)  (.O (in_int[508]), .I (in[438])) ;
    IBUF \in_ibuf(439)  (.O (in_int[509]), .I (in[439])) ;
    IBUF \in_ibuf(440)  (.O (in_int[510]), .I (in[440])) ;
    IBUF \in_ibuf(441)  (.O (in_int[511]), .I (in[441])) ;
    IBUF \in_ibuf(442)  (.O (in_int[512]), .I (in[442])) ;
    IBUF \in_ibuf(443)  (.O (in_int[513]), .I (in[443])) ;
    IBUF \in_ibuf(444)  (.O (in_int[514]), .I (in[444])) ;
    IBUF \in_ibuf(445)  (.O (in_int[515]), .I (in[445])) ;
    IBUF \in_ibuf(446)  (.O (in_int[516]), .I (in[446])) ;
    IBUF \in_ibuf(447)  (.O (in_int[517]), .I (in[447])) ;
    IBUF \in_ibuf(448)  (.O (in_int[518]), .I (in[448])) ;
    IBUF \in_ibuf(449)  (.O (in_int[519]), .I (in[449])) ;
    IBUF \in_ibuf(450)  (.O (in_int[520]), .I (in[450])) ;
    IBUF \in_ibuf(451)  (.O (in_int[521]), .I (in[451])) ;
    IBUF \in_ibuf(452)  (.O (in_int[522]), .I (in[452])) ;
    IBUF \in_ibuf(453)  (.O (in_int[523]), .I (in[453])) ;
    IBUF \in_ibuf(454)  (.O (in_int[524]), .I (in[454])) ;
    IBUF \in_ibuf(455)  (.O (in_int[525]), .I (in[455])) ;
    IBUF \in_ibuf(456)  (.O (in_int[526]), .I (in[456])) ;
    IBUF \in_ibuf(457)  (.O (in_int[527]), .I (in[457])) ;
    IBUF \in_ibuf(458)  (.O (in_int[528]), .I (in[458])) ;
    IBUF \in_ibuf(459)  (.O (in_int[529]), .I (in[459])) ;
    IBUF \in_ibuf(460)  (.O (in_int[530]), .I (in[460])) ;
    IBUF \in_ibuf(461)  (.O (in_int[531]), .I (in[461])) ;
    IBUF \in_ibuf(462)  (.O (in_int[532]), .I (in[462])) ;
    IBUF \in_ibuf(463)  (.O (in_int[533]), .I (in[463])) ;
    IBUF \in_ibuf(464)  (.O (in_int[534]), .I (in[464])) ;
    IBUF \in_ibuf(465)  (.O (in_int[535]), .I (in[465])) ;
    IBUF \in_ibuf(466)  (.O (in_int[536]), .I (in[466])) ;
    IBUF \in_ibuf(467)  (.O (in_int[537]), .I (in[467])) ;
    IBUF \in_ibuf(468)  (.O (in_int[538]), .I (in[468])) ;
    IBUF \in_ibuf(469)  (.O (in_int[539]), .I (in[469])) ;
    IBUF \in_ibuf(470)  (.O (in_int[540]), .I (in[470])) ;
    IBUF \in_ibuf(471)  (.O (in_int[541]), .I (in[471])) ;
    IBUF \in_ibuf(472)  (.O (in_int[542]), .I (in[472])) ;
    IBUF \in_ibuf(473)  (.O (in_int[543]), .I (in[473])) ;
    IBUF \in_ibuf(474)  (.O (in_int[544]), .I (in[474])) ;
    IBUF \in_ibuf(475)  (.O (in_int[545]), .I (in[475])) ;
    IBUF \in_ibuf(476)  (.O (in_int[546]), .I (in[476])) ;
    IBUF \in_ibuf(477)  (.O (in_int[547]), .I (in[477])) ;
    IBUF \in_ibuf(478)  (.O (in_int[548]), .I (in[478])) ;
    IBUF \in_ibuf(479)  (.O (in_int[549]), .I (in[479])) ;
    IBUF \in_ibuf(480)  (.O (in_int[550]), .I (in[480])) ;
    IBUF \in_ibuf(481)  (.O (in_int[551]), .I (in[481])) ;
    IBUF \in_ibuf(482)  (.O (in_int[552]), .I (in[482])) ;
    IBUF \in_ibuf(483)  (.O (in_int[553]), .I (in[483])) ;
    IBUF \in_ibuf(484)  (.O (in_int[554]), .I (in[484])) ;
    IBUF \in_ibuf(485)  (.O (in_int[555]), .I (in[485])) ;
    IBUF \in_ibuf(486)  (.O (in_int[556]), .I (in[486])) ;
    IBUF \in_ibuf(487)  (.O (in_int[557]), .I (in[487])) ;
    IBUF \in_ibuf(488)  (.O (in_int[558]), .I (in[488])) ;
    IBUF \in_ibuf(489)  (.O (in_int[559]), .I (in[489])) ;
    IBUF \in_ibuf(490)  (.O (in_int[560]), .I (in[490])) ;
    IBUF \in_ibuf(491)  (.O (in_int[561]), .I (in[491])) ;
    IBUF \in_ibuf(492)  (.O (in_int[562]), .I (in[492])) ;
    IBUF \in_ibuf(493)  (.O (in_int[563]), .I (in[493])) ;
    IBUF \in_ibuf(494)  (.O (in_int[564]), .I (in[494])) ;
    IBUF \in_ibuf(495)  (.O (in_int[565]), .I (in[495])) ;
    IBUF \in_ibuf(496)  (.O (in_int[566]), .I (in[496])) ;
    IBUF \in_ibuf(497)  (.O (in_int[567]), .I (in[497])) ;
    IBUF \in_ibuf(498)  (.O (in_int[568]), .I (in[498])) ;
    IBUF \in_ibuf(499)  (.O (in_int[569]), .I (in[499])) ;
    IBUF \in_ibuf(500)  (.O (in_int[570]), .I (in[500])) ;
    IBUF \in_ibuf(501)  (.O (in_int[571]), .I (in[501])) ;
    IBUF \in_ibuf(502)  (.O (in_int[572]), .I (in[502])) ;
    IBUF \in_ibuf(503)  (.O (in_int[573]), .I (in[503])) ;
    IBUF \in_ibuf(504)  (.O (in_int[574]), .I (in[504])) ;
    IBUF \in_ibuf(505)  (.O (in_int[575]), .I (in[505])) ;
    IBUF \in_ibuf(506)  (.O (in_int[576]), .I (in[506])) ;
    IBUF \in_ibuf(507)  (.O (in_int[577]), .I (in[507])) ;
    IBUF \in_ibuf(508)  (.O (in_int[578]), .I (in[508])) ;
    IBUF \in_ibuf(509)  (.O (in_int[579]), .I (in[509])) ;
    IBUF \in_ibuf(510)  (.O (in_int[580]), .I (in[510])) ;
    IBUF \in_ibuf(511)  (.O (in_int[581]), .I (in[511])) ;
    FD \reg_out(511)  (.Q (out_dup_0[511]), .D (in_int[70]), .C (clk_int)) ;
    FD \reg_out(510)  (.Q (out_dup_0[510]), .D (in_int[71]), .C (clk_int)) ;
    FD \reg_out(509)  (.Q (out_dup_0[509]), .D (in_int[72]), .C (clk_int)) ;
    FD \reg_out(508)  (.Q (out_dup_0[508]), .D (in_int[73]), .C (clk_int)) ;
    FD \reg_out(507)  (.Q (out_dup_0[507]), .D (in_int[74]), .C (clk_int)) ;
    FD \reg_out(506)  (.Q (out_dup_0[506]), .D (in_int[75]), .C (clk_int)) ;
    FD \reg_out(505)  (.Q (out_dup_0[505]), .D (in_int[76]), .C (clk_int)) ;
    FD \reg_out(504)  (.Q (out_dup_0[504]), .D (in_int[77]), .C (clk_int)) ;
    FD \reg_out(503)  (.Q (out_dup_0[503]), .D (in_int[78]), .C (clk_int)) ;
    FD \reg_out(502)  (.Q (out_dup_0[502]), .D (in_int[79]), .C (clk_int)) ;
    FD \reg_out(501)  (.Q (out_dup_0[501]), .D (in_int[80]), .C (clk_int)) ;
    FD \reg_out(500)  (.Q (out_dup_0[500]), .D (in_int[81]), .C (clk_int)) ;
    FD \reg_out(499)  (.Q (out_dup_0[499]), .D (in_int[82]), .C (clk_int)) ;
    FD \reg_out(498)  (.Q (out_dup_0[498]), .D (in_int[83]), .C (clk_int)) ;
    FD \reg_out(497)  (.Q (out_dup_0[497]), .D (in_int[84]), .C (clk_int)) ;
    FD \reg_out(496)  (.Q (out_dup_0[496]), .D (in_int[85]), .C (clk_int)) ;
    FD \reg_out(495)  (.Q (out_dup_0[495]), .D (in_int[86]), .C (clk_int)) ;
    FD \reg_out(494)  (.Q (out_dup_0[494]), .D (in_int[87]), .C (clk_int)) ;
    FD \reg_out(493)  (.Q (out_dup_0[493]), .D (in_int[88]), .C (clk_int)) ;
    FD \reg_out(492)  (.Q (out_dup_0[492]), .D (in_int[89]), .C (clk_int)) ;
    FD \reg_out(491)  (.Q (out_dup_0[491]), .D (in_int[90]), .C (clk_int)) ;
    FD \reg_out(490)  (.Q (out_dup_0[490]), .D (in_int[91]), .C (clk_int)) ;
    FD \reg_out(489)  (.Q (out_dup_0[489]), .D (in_int[92]), .C (clk_int)) ;
    FD \reg_out(488)  (.Q (out_dup_0[488]), .D (in_int[93]), .C (clk_int)) ;
    FD \reg_out(487)  (.Q (out_dup_0[487]), .D (in_int[94]), .C (clk_int)) ;
    FD \reg_out(486)  (.Q (out_dup_0[486]), .D (in_int[95]), .C (clk_int)) ;
    FD \reg_out(485)  (.Q (out_dup_0[485]), .D (in_int[96]), .C (clk_int)) ;
    FD \reg_out(484)  (.Q (out_dup_0[484]), .D (in_int[97]), .C (clk_int)) ;
    FD \reg_out(483)  (.Q (out_dup_0[483]), .D (in_int[98]), .C (clk_int)) ;
    FD \reg_out(482)  (.Q (out_dup_0[482]), .D (in_int[99]), .C (clk_int)) ;
    FD \reg_out(481)  (.Q (out_dup_0[481]), .D (in_int[100]), .C (clk_int)) ;
    FD \reg_out(480)  (.Q (out_dup_0[480]), .D (in_int[101]), .C (clk_int)) ;
    FD \reg_out(479)  (.Q (out_dup_0[479]), .D (in_int[102]), .C (clk_int)) ;
    FD \reg_out(478)  (.Q (out_dup_0[478]), .D (in_int[103]), .C (clk_int)) ;
    FD \reg_out(477)  (.Q (out_dup_0[477]), .D (in_int[104]), .C (clk_int)) ;
    FD \reg_out(476)  (.Q (out_dup_0[476]), .D (in_int[105]), .C (clk_int)) ;
    FD \reg_out(475)  (.Q (out_dup_0[475]), .D (in_int[106]), .C (clk_int)) ;
    FD \reg_out(474)  (.Q (out_dup_0[474]), .D (in_int[107]), .C (clk_int)) ;
    FD \reg_out(473)  (.Q (out_dup_0[473]), .D (in_int[108]), .C (clk_int)) ;
    FD \reg_out(472)  (.Q (out_dup_0[472]), .D (in_int[109]), .C (clk_int)) ;
    FD \reg_out(471)  (.Q (out_dup_0[471]), .D (in_int[110]), .C (clk_int)) ;
    FD \reg_out(470)  (.Q (out_dup_0[470]), .D (in_int[111]), .C (clk_int)) ;
    FD \reg_out(469)  (.Q (out_dup_0[469]), .D (in_int[112]), .C (clk_int)) ;
    FD \reg_out(468)  (.Q (out_dup_0[468]), .D (in_int[113]), .C (clk_int)) ;
    FD \reg_out(467)  (.Q (out_dup_0[467]), .D (in_int[114]), .C (clk_int)) ;
    FD \reg_out(466)  (.Q (out_dup_0[466]), .D (in_int[115]), .C (clk_int)) ;
    FD \reg_out(465)  (.Q (out_dup_0[465]), .D (in_int[116]), .C (clk_int)) ;
    FD \reg_out(464)  (.Q (out_dup_0[464]), .D (in_int[117]), .C (clk_int)) ;
    FD \reg_out(463)  (.Q (out_dup_0[463]), .D (in_int[118]), .C (clk_int)) ;
    FD \reg_out(462)  (.Q (out_dup_0[462]), .D (in_int[119]), .C (clk_int)) ;
    FD \reg_out(461)  (.Q (out_dup_0[461]), .D (in_int[120]), .C (clk_int)) ;
    FD \reg_out(460)  (.Q (out_dup_0[460]), .D (in_int[121]), .C (clk_int)) ;
    FD \reg_out(459)  (.Q (out_dup_0[459]), .D (in_int[122]), .C (clk_int)) ;
    FD \reg_out(458)  (.Q (out_dup_0[458]), .D (in_int[123]), .C (clk_int)) ;
    FD \reg_out(457)  (.Q (out_dup_0[457]), .D (in_int[124]), .C (clk_int)) ;
    FD \reg_out(456)  (.Q (out_dup_0[456]), .D (in_int[125]), .C (clk_int)) ;
    FD \reg_out(455)  (.Q (out_dup_0[455]), .D (in_int[126]), .C (clk_int)) ;
    FD \reg_out(454)  (.Q (out_dup_0[454]), .D (in_int[127]), .C (clk_int)) ;
    FD \reg_out(453)  (.Q (out_dup_0[453]), .D (in_int[128]), .C (clk_int)) ;
    FD \reg_out(452)  (.Q (out_dup_0[452]), .D (in_int[129]), .C (clk_int)) ;
    FD \reg_out(451)  (.Q (out_dup_0[451]), .D (in_int[130]), .C (clk_int)) ;
    FD \reg_out(450)  (.Q (out_dup_0[450]), .D (in_int[131]), .C (clk_int)) ;
    FD \reg_out(449)  (.Q (out_dup_0[449]), .D (in_int[132]), .C (clk_int)) ;
    FD \reg_out(448)  (.Q (out_dup_0[448]), .D (in_int[133]), .C (clk_int)) ;
    FD \reg_out(447)  (.Q (out_dup_0[447]), .D (in_int[134]), .C (clk_int)) ;
    FD \reg_out(446)  (.Q (out_dup_0[446]), .D (in_int[135]), .C (clk_int)) ;
    FD \reg_out(445)  (.Q (out_dup_0[445]), .D (in_int[136]), .C (clk_int)) ;
    FD \reg_out(444)  (.Q (out_dup_0[444]), .D (in_int[137]), .C (clk_int)) ;
    FD \reg_out(443)  (.Q (out_dup_0[443]), .D (in_int[138]), .C (clk_int)) ;
    FD \reg_out(442)  (.Q (out_dup_0[442]), .D (in_int[139]), .C (clk_int)) ;
    FD \reg_out(441)  (.Q (out_dup_0[441]), .D (in_int[140]), .C (clk_int)) ;
    FD \reg_out(440)  (.Q (out_dup_0[440]), .D (in_int[141]), .C (clk_int)) ;
    FD \reg_out(439)  (.Q (out_dup_0[439]), .D (in_int[142]), .C (clk_int)) ;
    FD \reg_out(438)  (.Q (out_dup_0[438]), .D (in_int[143]), .C (clk_int)) ;
    FD \reg_out(437)  (.Q (out_dup_0[437]), .D (in_int[144]), .C (clk_int)) ;
    FD \reg_out(436)  (.Q (out_dup_0[436]), .D (in_int[145]), .C (clk_int)) ;
    FD \reg_out(435)  (.Q (out_dup_0[435]), .D (in_int[146]), .C (clk_int)) ;
    FD \reg_out(434)  (.Q (out_dup_0[434]), .D (in_int[147]), .C (clk_int)) ;
    FD \reg_out(433)  (.Q (out_dup_0[433]), .D (in_int[148]), .C (clk_int)) ;
    FD \reg_out(432)  (.Q (out_dup_0[432]), .D (in_int[149]), .C (clk_int)) ;
    FD \reg_out(431)  (.Q (out_dup_0[431]), .D (in_int[150]), .C (clk_int)) ;
    FD \reg_out(430)  (.Q (out_dup_0[430]), .D (in_int[151]), .C (clk_int)) ;
    FD \reg_out(429)  (.Q (out_dup_0[429]), .D (in_int[152]), .C (clk_int)) ;
    FD \reg_out(428)  (.Q (out_dup_0[428]), .D (in_int[153]), .C (clk_int)) ;
    FD \reg_out(427)  (.Q (out_dup_0[427]), .D (in_int[154]), .C (clk_int)) ;
    FD \reg_out(426)  (.Q (out_dup_0[426]), .D (in_int[155]), .C (clk_int)) ;
    FD \reg_out(425)  (.Q (out_dup_0[425]), .D (in_int[156]), .C (clk_int)) ;
    FD \reg_out(424)  (.Q (out_dup_0[424]), .D (in_int[157]), .C (clk_int)) ;
    FD \reg_out(423)  (.Q (out_dup_0[423]), .D (in_int[158]), .C (clk_int)) ;
    FD \reg_out(422)  (.Q (out_dup_0[422]), .D (in_int[159]), .C (clk_int)) ;
    FD \reg_out(421)  (.Q (out_dup_0[421]), .D (in_int[160]), .C (clk_int)) ;
    FD \reg_out(420)  (.Q (out_dup_0[420]), .D (in_int[161]), .C (clk_int)) ;
    FD \reg_out(419)  (.Q (out_dup_0[419]), .D (in_int[162]), .C (clk_int)) ;
    FD \reg_out(418)  (.Q (out_dup_0[418]), .D (in_int[163]), .C (clk_int)) ;
    FD \reg_out(417)  (.Q (out_dup_0[417]), .D (in_int[164]), .C (clk_int)) ;
    FD \reg_out(416)  (.Q (out_dup_0[416]), .D (in_int[165]), .C (clk_int)) ;
    FD \reg_out(415)  (.Q (out_dup_0[415]), .D (in_int[166]), .C (clk_int)) ;
    FD \reg_out(414)  (.Q (out_dup_0[414]), .D (in_int[167]), .C (clk_int)) ;
    FD \reg_out(413)  (.Q (out_dup_0[413]), .D (in_int[168]), .C (clk_int)) ;
    FD \reg_out(412)  (.Q (out_dup_0[412]), .D (in_int[169]), .C (clk_int)) ;
    FD \reg_out(411)  (.Q (out_dup_0[411]), .D (in_int[170]), .C (clk_int)) ;
    FD \reg_out(410)  (.Q (out_dup_0[410]), .D (in_int[171]), .C (clk_int)) ;
    FD \reg_out(409)  (.Q (out_dup_0[409]), .D (in_int[172]), .C (clk_int)) ;
    FD \reg_out(408)  (.Q (out_dup_0[408]), .D (in_int[173]), .C (clk_int)) ;
    FD \reg_out(407)  (.Q (out_dup_0[407]), .D (in_int[174]), .C (clk_int)) ;
    FD \reg_out(406)  (.Q (out_dup_0[406]), .D (in_int[175]), .C (clk_int)) ;
    FD \reg_out(405)  (.Q (out_dup_0[405]), .D (in_int[176]), .C (clk_int)) ;
    FD \reg_out(404)  (.Q (out_dup_0[404]), .D (in_int[177]), .C (clk_int)) ;
    FD \reg_out(403)  (.Q (out_dup_0[403]), .D (in_int[178]), .C (clk_int)) ;
    FD \reg_out(402)  (.Q (out_dup_0[402]), .D (in_int[179]), .C (clk_int)) ;
    FD \reg_out(401)  (.Q (out_dup_0[401]), .D (in_int[180]), .C (clk_int)) ;
    FD \reg_out(400)  (.Q (out_dup_0[400]), .D (in_int[181]), .C (clk_int)) ;
    FD \reg_out(399)  (.Q (out_dup_0[399]), .D (in_int[182]), .C (clk_int)) ;
    FD \reg_out(398)  (.Q (out_dup_0[398]), .D (in_int[183]), .C (clk_int)) ;
    FD \reg_out(397)  (.Q (out_dup_0[397]), .D (in_int[184]), .C (clk_int)) ;
    FD \reg_out(396)  (.Q (out_dup_0[396]), .D (in_int[185]), .C (clk_int)) ;
    FD \reg_out(395)  (.Q (out_dup_0[395]), .D (in_int[186]), .C (clk_int)) ;
    FD \reg_out(394)  (.Q (out_dup_0[394]), .D (in_int[187]), .C (clk_int)) ;
    FD \reg_out(393)  (.Q (out_dup_0[393]), .D (in_int[188]), .C (clk_int)) ;
    FD \reg_out(392)  (.Q (out_dup_0[392]), .D (in_int[189]), .C (clk_int)) ;
    FD \reg_out(391)  (.Q (out_dup_0[391]), .D (in_int[190]), .C (clk_int)) ;
    FD \reg_out(390)  (.Q (out_dup_0[390]), .D (in_int[191]), .C (clk_int)) ;
    FD \reg_out(389)  (.Q (out_dup_0[389]), .D (in_int[192]), .C (clk_int)) ;
    FD \reg_out(388)  (.Q (out_dup_0[388]), .D (in_int[193]), .C (clk_int)) ;
    FD \reg_out(387)  (.Q (out_dup_0[387]), .D (in_int[194]), .C (clk_int)) ;
    FD \reg_out(386)  (.Q (out_dup_0[386]), .D (in_int[195]), .C (clk_int)) ;
    FD \reg_out(385)  (.Q (out_dup_0[385]), .D (in_int[196]), .C (clk_int)) ;
    FD \reg_out(384)  (.Q (out_dup_0[384]), .D (in_int[197]), .C (clk_int)) ;
    FD \reg_out(383)  (.Q (out_dup_0[383]), .D (in_int[198]), .C (clk_int)) ;
    FD \reg_out(382)  (.Q (out_dup_0[382]), .D (in_int[199]), .C (clk_int)) ;
    FD \reg_out(381)  (.Q (out_dup_0[381]), .D (in_int[200]), .C (clk_int)) ;
    FD \reg_out(380)  (.Q (out_dup_0[380]), .D (in_int[201]), .C (clk_int)) ;
    FD \reg_out(379)  (.Q (out_dup_0[379]), .D (in_int[202]), .C (clk_int)) ;
    FD \reg_out(378)  (.Q (out_dup_0[378]), .D (in_int[203]), .C (clk_int)) ;
    FD \reg_out(377)  (.Q (out_dup_0[377]), .D (in_int[204]), .C (clk_int)) ;
    FD \reg_out(376)  (.Q (out_dup_0[376]), .D (in_int[205]), .C (clk_int)) ;
    FD \reg_out(375)  (.Q (out_dup_0[375]), .D (in_int[206]), .C (clk_int)) ;
    FD \reg_out(374)  (.Q (out_dup_0[374]), .D (in_int[207]), .C (clk_int)) ;
    FD \reg_out(373)  (.Q (out_dup_0[373]), .D (in_int[208]), .C (clk_int)) ;
    FD \reg_out(372)  (.Q (out_dup_0[372]), .D (in_int[209]), .C (clk_int)) ;
    FD \reg_out(371)  (.Q (out_dup_0[371]), .D (in_int[210]), .C (clk_int)) ;
    FD \reg_out(370)  (.Q (out_dup_0[370]), .D (in_int[211]), .C (clk_int)) ;
    FD \reg_out(369)  (.Q (out_dup_0[369]), .D (in_int[212]), .C (clk_int)) ;
    FD \reg_out(368)  (.Q (out_dup_0[368]), .D (in_int[213]), .C (clk_int)) ;
    FD \reg_out(367)  (.Q (out_dup_0[367]), .D (in_int[214]), .C (clk_int)) ;
    FD \reg_out(366)  (.Q (out_dup_0[366]), .D (in_int[215]), .C (clk_int)) ;
    FD \reg_out(365)  (.Q (out_dup_0[365]), .D (in_int[216]), .C (clk_int)) ;
    FD \reg_out(364)  (.Q (out_dup_0[364]), .D (in_int[217]), .C (clk_int)) ;
    FD \reg_out(363)  (.Q (out_dup_0[363]), .D (in_int[218]), .C (clk_int)) ;
    FD \reg_out(362)  (.Q (out_dup_0[362]), .D (in_int[219]), .C (clk_int)) ;
    FD \reg_out(361)  (.Q (out_dup_0[361]), .D (in_int[220]), .C (clk_int)) ;
    FD \reg_out(360)  (.Q (out_dup_0[360]), .D (in_int[221]), .C (clk_int)) ;
    FD \reg_out(359)  (.Q (out_dup_0[359]), .D (in_int[222]), .C (clk_int)) ;
    FD \reg_out(358)  (.Q (out_dup_0[358]), .D (in_int[223]), .C (clk_int)) ;
    FD \reg_out(357)  (.Q (out_dup_0[357]), .D (in_int[224]), .C (clk_int)) ;
    FD \reg_out(356)  (.Q (out_dup_0[356]), .D (in_int[225]), .C (clk_int)) ;
    FD \reg_out(355)  (.Q (out_dup_0[355]), .D (in_int[226]), .C (clk_int)) ;
    FD \reg_out(354)  (.Q (out_dup_0[354]), .D (in_int[227]), .C (clk_int)) ;
    FD \reg_out(353)  (.Q (out_dup_0[353]), .D (in_int[228]), .C (clk_int)) ;
    FD \reg_out(352)  (.Q (out_dup_0[352]), .D (in_int[229]), .C (clk_int)) ;
    FD \reg_out(351)  (.Q (out_dup_0[351]), .D (in_int[230]), .C (clk_int)) ;
    FD \reg_out(350)  (.Q (out_dup_0[350]), .D (in_int[231]), .C (clk_int)) ;
    FD \reg_out(349)  (.Q (out_dup_0[349]), .D (in_int[232]), .C (clk_int)) ;
    FD \reg_out(348)  (.Q (out_dup_0[348]), .D (in_int[233]), .C (clk_int)) ;
    FD \reg_out(347)  (.Q (out_dup_0[347]), .D (in_int[234]), .C (clk_int)) ;
    FD \reg_out(346)  (.Q (out_dup_0[346]), .D (in_int[235]), .C (clk_int)) ;
    FD \reg_out(345)  (.Q (out_dup_0[345]), .D (in_int[236]), .C (clk_int)) ;
    FD \reg_out(344)  (.Q (out_dup_0[344]), .D (in_int[237]), .C (clk_int)) ;
    FD \reg_out(343)  (.Q (out_dup_0[343]), .D (in_int[238]), .C (clk_int)) ;
    FD \reg_out(342)  (.Q (out_dup_0[342]), .D (in_int[239]), .C (clk_int)) ;
    FD \reg_out(341)  (.Q (out_dup_0[341]), .D (in_int[240]), .C (clk_int)) ;
    FD \reg_out(340)  (.Q (out_dup_0[340]), .D (in_int[241]), .C (clk_int)) ;
    FD \reg_out(339)  (.Q (out_dup_0[339]), .D (in_int[242]), .C (clk_int)) ;
    FD \reg_out(338)  (.Q (out_dup_0[338]), .D (in_int[243]), .C (clk_int)) ;
    FD \reg_out(337)  (.Q (out_dup_0[337]), .D (in_int[244]), .C (clk_int)) ;
    FD \reg_out(336)  (.Q (out_dup_0[336]), .D (in_int[245]), .C (clk_int)) ;
    FD \reg_out(335)  (.Q (out_dup_0[335]), .D (in_int[246]), .C (clk_int)) ;
    FD \reg_out(334)  (.Q (out_dup_0[334]), .D (in_int[247]), .C (clk_int)) ;
    FD \reg_out(333)  (.Q (out_dup_0[333]), .D (in_int[248]), .C (clk_int)) ;
    FD \reg_out(332)  (.Q (out_dup_0[332]), .D (in_int[249]), .C (clk_int)) ;
    FD \reg_out(331)  (.Q (out_dup_0[331]), .D (in_int[250]), .C (clk_int)) ;
    FD \reg_out(330)  (.Q (out_dup_0[330]), .D (in_int[251]), .C (clk_int)) ;
    FD \reg_out(329)  (.Q (out_dup_0[329]), .D (in_int[252]), .C (clk_int)) ;
    FD \reg_out(328)  (.Q (out_dup_0[328]), .D (in_int[253]), .C (clk_int)) ;
    FD \reg_out(327)  (.Q (out_dup_0[327]), .D (in_int[254]), .C (clk_int)) ;
    FD \reg_out(326)  (.Q (out_dup_0[326]), .D (in_int[255]), .C (clk_int)) ;
    FD \reg_out(325)  (.Q (out_dup_0[325]), .D (in_int[256]), .C (clk_int)) ;
    FD \reg_out(324)  (.Q (out_dup_0[324]), .D (in_int[257]), .C (clk_int)) ;
    FD \reg_out(323)  (.Q (out_dup_0[323]), .D (in_int[258]), .C (clk_int)) ;
    FD \reg_out(322)  (.Q (out_dup_0[322]), .D (in_int[259]), .C (clk_int)) ;
    FD \reg_out(321)  (.Q (out_dup_0[321]), .D (in_int[260]), .C (clk_int)) ;
    FD \reg_out(320)  (.Q (out_dup_0[320]), .D (in_int[261]), .C (clk_int)) ;
    FD \reg_out(319)  (.Q (out_dup_0[319]), .D (in_int[262]), .C (clk_int)) ;
    FD \reg_out(318)  (.Q (out_dup_0[318]), .D (in_int[263]), .C (clk_int)) ;
    FD \reg_out(317)  (.Q (out_dup_0[317]), .D (in_int[264]), .C (clk_int)) ;
    FD \reg_out(316)  (.Q (out_dup_0[316]), .D (in_int[265]), .C (clk_int)) ;
    FD \reg_out(315)  (.Q (out_dup_0[315]), .D (in_int[266]), .C (clk_int)) ;
    FD \reg_out(314)  (.Q (out_dup_0[314]), .D (in_int[267]), .C (clk_int)) ;
    FD \reg_out(313)  (.Q (out_dup_0[313]), .D (in_int[268]), .C (clk_int)) ;
    FD \reg_out(312)  (.Q (out_dup_0[312]), .D (in_int[269]), .C (clk_int)) ;
    FD \reg_out(311)  (.Q (out_dup_0[311]), .D (in_int[270]), .C (clk_int)) ;
    FD \reg_out(310)  (.Q (out_dup_0[310]), .D (in_int[271]), .C (clk_int)) ;
    FD \reg_out(309)  (.Q (out_dup_0[309]), .D (in_int[272]), .C (clk_int)) ;
    FD \reg_out(308)  (.Q (out_dup_0[308]), .D (in_int[273]), .C (clk_int)) ;
    FD \reg_out(307)  (.Q (out_dup_0[307]), .D (in_int[274]), .C (clk_int)) ;
    FD \reg_out(306)  (.Q (out_dup_0[306]), .D (in_int[275]), .C (clk_int)) ;
    FD \reg_out(305)  (.Q (out_dup_0[305]), .D (in_int[276]), .C (clk_int)) ;
    FD \reg_out(304)  (.Q (out_dup_0[304]), .D (in_int[277]), .C (clk_int)) ;
    FD \reg_out(303)  (.Q (out_dup_0[303]), .D (in_int[278]), .C (clk_int)) ;
    FD \reg_out(302)  (.Q (out_dup_0[302]), .D (in_int[279]), .C (clk_int)) ;
    FD \reg_out(301)  (.Q (out_dup_0[301]), .D (in_int[280]), .C (clk_int)) ;
    FD \reg_out(300)  (.Q (out_dup_0[300]), .D (in_int[281]), .C (clk_int)) ;
    FD \reg_out(299)  (.Q (out_dup_0[299]), .D (in_int[282]), .C (clk_int)) ;
    FD \reg_out(298)  (.Q (out_dup_0[298]), .D (in_int[283]), .C (clk_int)) ;
    FD \reg_out(297)  (.Q (out_dup_0[297]), .D (in_int[284]), .C (clk_int)) ;
    FD \reg_out(296)  (.Q (out_dup_0[296]), .D (in_int[285]), .C (clk_int)) ;
    FD \reg_out(295)  (.Q (out_dup_0[295]), .D (in_int[286]), .C (clk_int)) ;
    FD \reg_out(294)  (.Q (out_dup_0[294]), .D (in_int[287]), .C (clk_int)) ;
    FD \reg_out(293)  (.Q (out_dup_0[293]), .D (in_int[288]), .C (clk_int)) ;
    FD \reg_out(292)  (.Q (out_dup_0[292]), .D (in_int[289]), .C (clk_int)) ;
    FD \reg_out(291)  (.Q (out_dup_0[291]), .D (in_int[290]), .C (clk_int)) ;
    FD \reg_out(290)  (.Q (out_dup_0[290]), .D (in_int[291]), .C (clk_int)) ;
    FD \reg_out(289)  (.Q (out_dup_0[289]), .D (in_int[292]), .C (clk_int)) ;
    FD \reg_out(288)  (.Q (out_dup_0[288]), .D (in_int[293]), .C (clk_int)) ;
    FD \reg_out(287)  (.Q (out_dup_0[287]), .D (in_int[294]), .C (clk_int)) ;
    FD \reg_out(286)  (.Q (out_dup_0[286]), .D (in_int[295]), .C (clk_int)) ;
    FD \reg_out(285)  (.Q (out_dup_0[285]), .D (in_int[296]), .C (clk_int)) ;
    FD \reg_out(284)  (.Q (out_dup_0[284]), .D (in_int[297]), .C (clk_int)) ;
    FD \reg_out(283)  (.Q (out_dup_0[283]), .D (in_int[298]), .C (clk_int)) ;
    FD \reg_out(282)  (.Q (out_dup_0[282]), .D (in_int[299]), .C (clk_int)) ;
    FD \reg_out(281)  (.Q (out_dup_0[281]), .D (in_int[300]), .C (clk_int)) ;
    FD \reg_out(280)  (.Q (out_dup_0[280]), .D (in_int[301]), .C (clk_int)) ;
    FD \reg_out(279)  (.Q (out_dup_0[279]), .D (in_int[302]), .C (clk_int)) ;
    FD \reg_out(278)  (.Q (out_dup_0[278]), .D (in_int[303]), .C (clk_int)) ;
    FD \reg_out(277)  (.Q (out_dup_0[277]), .D (in_int[304]), .C (clk_int)) ;
    FD \reg_out(276)  (.Q (out_dup_0[276]), .D (in_int[305]), .C (clk_int)) ;
    FD \reg_out(275)  (.Q (out_dup_0[275]), .D (in_int[306]), .C (clk_int)) ;
    FD \reg_out(274)  (.Q (out_dup_0[274]), .D (in_int[307]), .C (clk_int)) ;
    FD \reg_out(273)  (.Q (out_dup_0[273]), .D (in_int[308]), .C (clk_int)) ;
    FD \reg_out(272)  (.Q (out_dup_0[272]), .D (in_int[309]), .C (clk_int)) ;
    FD \reg_out(271)  (.Q (out_dup_0[271]), .D (in_int[310]), .C (clk_int)) ;
    FD \reg_out(270)  (.Q (out_dup_0[270]), .D (in_int[311]), .C (clk_int)) ;
    FD \reg_out(269)  (.Q (out_dup_0[269]), .D (in_int[312]), .C (clk_int)) ;
    FD \reg_out(268)  (.Q (out_dup_0[268]), .D (in_int[313]), .C (clk_int)) ;
    FD \reg_out(267)  (.Q (out_dup_0[267]), .D (in_int[314]), .C (clk_int)) ;
    FD \reg_out(266)  (.Q (out_dup_0[266]), .D (in_int[315]), .C (clk_int)) ;
    FD \reg_out(265)  (.Q (out_dup_0[265]), .D (in_int[316]), .C (clk_int)) ;
    FD \reg_out(264)  (.Q (out_dup_0[264]), .D (in_int[317]), .C (clk_int)) ;
    FD \reg_out(263)  (.Q (out_dup_0[263]), .D (in_int[318]), .C (clk_int)) ;
    FD \reg_out(262)  (.Q (out_dup_0[262]), .D (in_int[319]), .C (clk_int)) ;
    FD \reg_out(261)  (.Q (out_dup_0[261]), .D (in_int[320]), .C (clk_int)) ;
    FD \reg_out(260)  (.Q (out_dup_0[260]), .D (in_int[321]), .C (clk_int)) ;
    FD \reg_out(259)  (.Q (out_dup_0[259]), .D (in_int[322]), .C (clk_int)) ;
    FD \reg_out(258)  (.Q (out_dup_0[258]), .D (in_int[323]), .C (clk_int)) ;
    FD \reg_out(257)  (.Q (out_dup_0[257]), .D (in_int[324]), .C (clk_int)) ;
    FD \reg_out(256)  (.Q (out_dup_0[256]), .D (in_int[325]), .C (clk_int)) ;
    FD \reg_out(255)  (.Q (out_dup_0[255]), .D (in_int[326]), .C (clk_int)) ;
    FD \reg_out(254)  (.Q (out_dup_0[254]), .D (in_int[327]), .C (clk_int)) ;
    FD \reg_out(253)  (.Q (out_dup_0[253]), .D (in_int[328]), .C (clk_int)) ;
    FD \reg_out(252)  (.Q (out_dup_0[252]), .D (in_int[329]), .C (clk_int)) ;
    FD \reg_out(251)  (.Q (out_dup_0[251]), .D (in_int[330]), .C (clk_int)) ;
    FD \reg_out(250)  (.Q (out_dup_0[250]), .D (in_int[331]), .C (clk_int)) ;
    FD \reg_out(249)  (.Q (out_dup_0[249]), .D (in_int[332]), .C (clk_int)) ;
    FD \reg_out(248)  (.Q (out_dup_0[248]), .D (in_int[333]), .C (clk_int)) ;
    FD \reg_out(247)  (.Q (out_dup_0[247]), .D (in_int[334]), .C (clk_int)) ;
    FD \reg_out(246)  (.Q (out_dup_0[246]), .D (in_int[335]), .C (clk_int)) ;
    FD \reg_out(245)  (.Q (out_dup_0[245]), .D (in_int[336]), .C (clk_int)) ;
    FD \reg_out(244)  (.Q (out_dup_0[244]), .D (in_int[337]), .C (clk_int)) ;
    FD \reg_out(243)  (.Q (out_dup_0[243]), .D (in_int[338]), .C (clk_int)) ;
    FD \reg_out(242)  (.Q (out_dup_0[242]), .D (in_int[339]), .C (clk_int)) ;
    FD \reg_out(241)  (.Q (out_dup_0[241]), .D (in_int[340]), .C (clk_int)) ;
    FD \reg_out(240)  (.Q (out_dup_0[240]), .D (in_int[341]), .C (clk_int)) ;
    FD \reg_out(239)  (.Q (out_dup_0[239]), .D (in_int[342]), .C (clk_int)) ;
    FD \reg_out(238)  (.Q (out_dup_0[238]), .D (in_int[343]), .C (clk_int)) ;
    FD \reg_out(237)  (.Q (out_dup_0[237]), .D (in_int[344]), .C (clk_int)) ;
    FD \reg_out(236)  (.Q (out_dup_0[236]), .D (in_int[345]), .C (clk_int)) ;
    FD \reg_out(235)  (.Q (out_dup_0[235]), .D (in_int[346]), .C (clk_int)) ;
    FD \reg_out(234)  (.Q (out_dup_0[234]), .D (in_int[347]), .C (clk_int)) ;
    FD \reg_out(233)  (.Q (out_dup_0[233]), .D (in_int[348]), .C (clk_int)) ;
    FD \reg_out(232)  (.Q (out_dup_0[232]), .D (in_int[349]), .C (clk_int)) ;
    FD \reg_out(231)  (.Q (out_dup_0[231]), .D (in_int[350]), .C (clk_int)) ;
    FD \reg_out(230)  (.Q (out_dup_0[230]), .D (in_int[351]), .C (clk_int)) ;
    FD \reg_out(229)  (.Q (out_dup_0[229]), .D (in_int[352]), .C (clk_int)) ;
    FD \reg_out(228)  (.Q (out_dup_0[228]), .D (in_int[353]), .C (clk_int)) ;
    FD \reg_out(227)  (.Q (out_dup_0[227]), .D (in_int[354]), .C (clk_int)) ;
    FD \reg_out(226)  (.Q (out_dup_0[226]), .D (in_int[355]), .C (clk_int)) ;
    FD \reg_out(225)  (.Q (out_dup_0[225]), .D (in_int[356]), .C (clk_int)) ;
    FD \reg_out(224)  (.Q (out_dup_0[224]), .D (in_int[357]), .C (clk_int)) ;
    FD \reg_out(223)  (.Q (out_dup_0[223]), .D (in_int[358]), .C (clk_int)) ;
    FD \reg_out(222)  (.Q (out_dup_0[222]), .D (in_int[359]), .C (clk_int)) ;
    FD \reg_out(221)  (.Q (out_dup_0[221]), .D (in_int[360]), .C (clk_int)) ;
    FD \reg_out(220)  (.Q (out_dup_0[220]), .D (in_int[361]), .C (clk_int)) ;
    FD \reg_out(219)  (.Q (out_dup_0[219]), .D (in_int[362]), .C (clk_int)) ;
    FD \reg_out(218)  (.Q (out_dup_0[218]), .D (in_int[363]), .C (clk_int)) ;
    FD \reg_out(217)  (.Q (out_dup_0[217]), .D (in_int[364]), .C (clk_int)) ;
    FD \reg_out(216)  (.Q (out_dup_0[216]), .D (in_int[365]), .C (clk_int)) ;
    FD \reg_out(215)  (.Q (out_dup_0[215]), .D (in_int[366]), .C (clk_int)) ;
    FD \reg_out(214)  (.Q (out_dup_0[214]), .D (in_int[367]), .C (clk_int)) ;
    FD \reg_out(213)  (.Q (out_dup_0[213]), .D (in_int[368]), .C (clk_int)) ;
    FD \reg_out(212)  (.Q (out_dup_0[212]), .D (in_int[369]), .C (clk_int)) ;
    FD \reg_out(211)  (.Q (out_dup_0[211]), .D (in_int[370]), .C (clk_int)) ;
    FD \reg_out(210)  (.Q (out_dup_0[210]), .D (in_int[371]), .C (clk_int)) ;
    FD \reg_out(209)  (.Q (out_dup_0[209]), .D (in_int[372]), .C (clk_int)) ;
    FD \reg_out(208)  (.Q (out_dup_0[208]), .D (in_int[373]), .C (clk_int)) ;
    FD \reg_out(207)  (.Q (out_dup_0[207]), .D (in_int[374]), .C (clk_int)) ;
    FD \reg_out(206)  (.Q (out_dup_0[206]), .D (in_int[375]), .C (clk_int)) ;
    FD \reg_out(205)  (.Q (out_dup_0[205]), .D (in_int[376]), .C (clk_int)) ;
    FD \reg_out(204)  (.Q (out_dup_0[204]), .D (in_int[377]), .C (clk_int)) ;
    FD \reg_out(203)  (.Q (out_dup_0[203]), .D (in_int[378]), .C (clk_int)) ;
    FD \reg_out(202)  (.Q (out_dup_0[202]), .D (in_int[379]), .C (clk_int)) ;
    FD \reg_out(201)  (.Q (out_dup_0[201]), .D (in_int[380]), .C (clk_int)) ;
    FD \reg_out(200)  (.Q (out_dup_0[200]), .D (in_int[381]), .C (clk_int)) ;
    FD \reg_out(199)  (.Q (out_dup_0[199]), .D (in_int[382]), .C (clk_int)) ;
    FD \reg_out(198)  (.Q (out_dup_0[198]), .D (in_int[383]), .C (clk_int)) ;
    FD \reg_out(197)  (.Q (out_dup_0[197]), .D (in_int[384]), .C (clk_int)) ;
    FD \reg_out(196)  (.Q (out_dup_0[196]), .D (in_int[385]), .C (clk_int)) ;
    FD \reg_out(195)  (.Q (out_dup_0[195]), .D (in_int[386]), .C (clk_int)) ;
    FD \reg_out(194)  (.Q (out_dup_0[194]), .D (in_int[387]), .C (clk_int)) ;
    FD \reg_out(193)  (.Q (out_dup_0[193]), .D (in_int[388]), .C (clk_int)) ;
    FD \reg_out(192)  (.Q (out_dup_0[192]), .D (in_int[389]), .C (clk_int)) ;
    FD \reg_out(191)  (.Q (out_dup_0[191]), .D (in_int[390]), .C (clk_int)) ;
    FD \reg_out(190)  (.Q (out_dup_0[190]), .D (in_int[391]), .C (clk_int)) ;
    FD \reg_out(189)  (.Q (out_dup_0[189]), .D (in_int[392]), .C (clk_int)) ;
    FD \reg_out(188)  (.Q (out_dup_0[188]), .D (in_int[393]), .C (clk_int)) ;
    FD \reg_out(187)  (.Q (out_dup_0[187]), .D (in_int[394]), .C (clk_int)) ;
    FD \reg_out(186)  (.Q (out_dup_0[186]), .D (in_int[395]), .C (clk_int)) ;
    FD \reg_out(185)  (.Q (out_dup_0[185]), .D (in_int[396]), .C (clk_int)) ;
    FD \reg_out(184)  (.Q (out_dup_0[184]), .D (in_int[397]), .C (clk_int)) ;
    FD \reg_out(183)  (.Q (out_dup_0[183]), .D (in_int[398]), .C (clk_int)) ;
    FD \reg_out(182)  (.Q (out_dup_0[182]), .D (in_int[399]), .C (clk_int)) ;
    FD \reg_out(181)  (.Q (out_dup_0[181]), .D (in_int[400]), .C (clk_int)) ;
    FD \reg_out(180)  (.Q (out_dup_0[180]), .D (in_int[401]), .C (clk_int)) ;
    FD \reg_out(179)  (.Q (out_dup_0[179]), .D (in_int[402]), .C (clk_int)) ;
    FD \reg_out(178)  (.Q (out_dup_0[178]), .D (in_int[403]), .C (clk_int)) ;
    FD \reg_out(177)  (.Q (out_dup_0[177]), .D (in_int[404]), .C (clk_int)) ;
    FD \reg_out(176)  (.Q (out_dup_0[176]), .D (in_int[405]), .C (clk_int)) ;
    FD \reg_out(175)  (.Q (out_dup_0[175]), .D (in_int[406]), .C (clk_int)) ;
    FD \reg_out(174)  (.Q (out_dup_0[174]), .D (in_int[407]), .C (clk_int)) ;
    FD \reg_out(173)  (.Q (out_dup_0[173]), .D (in_int[408]), .C (clk_int)) ;
    FD \reg_out(172)  (.Q (out_dup_0[172]), .D (in_int[409]), .C (clk_int)) ;
    FD \reg_out(171)  (.Q (out_dup_0[171]), .D (in_int[410]), .C (clk_int)) ;
    FD \reg_out(170)  (.Q (out_dup_0[170]), .D (in_int[411]), .C (clk_int)) ;
    FD \reg_out(169)  (.Q (out_dup_0[169]), .D (in_int[412]), .C (clk_int)) ;
    FD \reg_out(168)  (.Q (out_dup_0[168]), .D (in_int[413]), .C (clk_int)) ;
    FD \reg_out(167)  (.Q (out_dup_0[167]), .D (in_int[414]), .C (clk_int)) ;
    FD \reg_out(166)  (.Q (out_dup_0[166]), .D (in_int[415]), .C (clk_int)) ;
    FD \reg_out(165)  (.Q (out_dup_0[165]), .D (in_int[416]), .C (clk_int)) ;
    FD \reg_out(164)  (.Q (out_dup_0[164]), .D (in_int[417]), .C (clk_int)) ;
    FD \reg_out(163)  (.Q (out_dup_0[163]), .D (in_int[418]), .C (clk_int)) ;
    FD \reg_out(162)  (.Q (out_dup_0[162]), .D (in_int[419]), .C (clk_int)) ;
    FD \reg_out(161)  (.Q (out_dup_0[161]), .D (in_int[420]), .C (clk_int)) ;
    FD \reg_out(160)  (.Q (out_dup_0[160]), .D (in_int[421]), .C (clk_int)) ;
    FD \reg_out(159)  (.Q (out_dup_0[159]), .D (in_int[422]), .C (clk_int)) ;
    FD \reg_out(158)  (.Q (out_dup_0[158]), .D (in_int[423]), .C (clk_int)) ;
    FD \reg_out(157)  (.Q (out_dup_0[157]), .D (in_int[424]), .C (clk_int)) ;
    FD \reg_out(156)  (.Q (out_dup_0[156]), .D (in_int[425]), .C (clk_int)) ;
    FD \reg_out(155)  (.Q (out_dup_0[155]), .D (in_int[426]), .C (clk_int)) ;
    FD \reg_out(154)  (.Q (out_dup_0[154]), .D (in_int[427]), .C (clk_int)) ;
    FD \reg_out(153)  (.Q (out_dup_0[153]), .D (in_int[428]), .C (clk_int)) ;
    FD \reg_out(152)  (.Q (out_dup_0[152]), .D (in_int[429]), .C (clk_int)) ;
    FD \reg_out(151)  (.Q (out_dup_0[151]), .D (in_int[430]), .C (clk_int)) ;
    FD \reg_out(150)  (.Q (out_dup_0[150]), .D (in_int[431]), .C (clk_int)) ;
    FD \reg_out(149)  (.Q (out_dup_0[149]), .D (in_int[432]), .C (clk_int)) ;
    FD \reg_out(148)  (.Q (out_dup_0[148]), .D (in_int[433]), .C (clk_int)) ;
    FD \reg_out(147)  (.Q (out_dup_0[147]), .D (in_int[434]), .C (clk_int)) ;
    FD \reg_out(146)  (.Q (out_dup_0[146]), .D (in_int[435]), .C (clk_int)) ;
    FD \reg_out(145)  (.Q (out_dup_0[145]), .D (in_int[436]), .C (clk_int)) ;
    FD \reg_out(144)  (.Q (out_dup_0[144]), .D (in_int[437]), .C (clk_int)) ;
    FD \reg_out(143)  (.Q (out_dup_0[143]), .D (in_int[438]), .C (clk_int)) ;
    FD \reg_out(142)  (.Q (out_dup_0[142]), .D (in_int[439]), .C (clk_int)) ;
    FD \reg_out(141)  (.Q (out_dup_0[141]), .D (in_int[440]), .C (clk_int)) ;
    FD \reg_out(140)  (.Q (out_dup_0[140]), .D (in_int[441]), .C (clk_int)) ;
    FD \reg_out(139)  (.Q (out_dup_0[139]), .D (in_int[442]), .C (clk_int)) ;
    FD \reg_out(138)  (.Q (out_dup_0[138]), .D (in_int[443]), .C (clk_int)) ;
    FD \reg_out(137)  (.Q (out_dup_0[137]), .D (in_int[444]), .C (clk_int)) ;
    FD \reg_out(136)  (.Q (out_dup_0[136]), .D (in_int[445]), .C (clk_int)) ;
    FD \reg_out(135)  (.Q (out_dup_0[135]), .D (in_int[446]), .C (clk_int)) ;
    FD \reg_out(134)  (.Q (out_dup_0[134]), .D (in_int[447]), .C (clk_int)) ;
    FD \reg_out(133)  (.Q (out_dup_0[133]), .D (in_int[448]), .C (clk_int)) ;
    FD \reg_out(132)  (.Q (out_dup_0[132]), .D (in_int[449]), .C (clk_int)) ;
    FD \reg_out(131)  (.Q (out_dup_0[131]), .D (in_int[450]), .C (clk_int)) ;
    FD \reg_out(130)  (.Q (out_dup_0[130]), .D (in_int[451]), .C (clk_int)) ;
    FD \reg_out(129)  (.Q (out_dup_0[129]), .D (in_int[452]), .C (clk_int)) ;
    FD \reg_out(128)  (.Q (out_dup_0[128]), .D (in_int[453]), .C (clk_int)) ;
    FD \reg_out(127)  (.Q (out_dup_0[127]), .D (in_int[454]), .C (clk_int)) ;
    FD \reg_out(126)  (.Q (out_dup_0[126]), .D (in_int[455]), .C (clk_int)) ;
    FD \reg_out(125)  (.Q (out_dup_0[125]), .D (in_int[456]), .C (clk_int)) ;
    FD \reg_out(124)  (.Q (out_dup_0[124]), .D (in_int[457]), .C (clk_int)) ;
    FD \reg_out(123)  (.Q (out_dup_0[123]), .D (in_int[458]), .C (clk_int)) ;
    FD \reg_out(122)  (.Q (out_dup_0[122]), .D (in_int[459]), .C (clk_int)) ;
    FD \reg_out(121)  (.Q (out_dup_0[121]), .D (in_int[460]), .C (clk_int)) ;
    FD \reg_out(120)  (.Q (out_dup_0[120]), .D (in_int[461]), .C (clk_int)) ;
    FD \reg_out(119)  (.Q (out_dup_0[119]), .D (in_int[462]), .C (clk_int)) ;
    FD \reg_out(118)  (.Q (out_dup_0[118]), .D (in_int[463]), .C (clk_int)) ;
    FD \reg_out(117)  (.Q (out_dup_0[117]), .D (in_int[464]), .C (clk_int)) ;
    FD \reg_out(116)  (.Q (out_dup_0[116]), .D (in_int[465]), .C (clk_int)) ;
    FD \reg_out(115)  (.Q (out_dup_0[115]), .D (in_int[466]), .C (clk_int)) ;
    FD \reg_out(114)  (.Q (out_dup_0[114]), .D (in_int[467]), .C (clk_int)) ;
    FD \reg_out(113)  (.Q (out_dup_0[113]), .D (in_int[468]), .C (clk_int)) ;
    FD \reg_out(112)  (.Q (out_dup_0[112]), .D (in_int[469]), .C (clk_int)) ;
    FD \reg_out(111)  (.Q (out_dup_0[111]), .D (in_int[470]), .C (clk_int)) ;
    FD \reg_out(110)  (.Q (out_dup_0[110]), .D (in_int[471]), .C (clk_int)) ;
    FD \reg_out(109)  (.Q (out_dup_0[109]), .D (in_int[472]), .C (clk_int)) ;
    FD \reg_out(108)  (.Q (out_dup_0[108]), .D (in_int[473]), .C (clk_int)) ;
    FD \reg_out(107)  (.Q (out_dup_0[107]), .D (in_int[474]), .C (clk_int)) ;
    FD \reg_out(106)  (.Q (out_dup_0[106]), .D (in_int[475]), .C (clk_int)) ;
    FD \reg_out(105)  (.Q (out_dup_0[105]), .D (in_int[476]), .C (clk_int)) ;
    FD \reg_out(104)  (.Q (out_dup_0[104]), .D (in_int[477]), .C (clk_int)) ;
    FD \reg_out(103)  (.Q (out_dup_0[103]), .D (in_int[478]), .C (clk_int)) ;
    FD \reg_out(102)  (.Q (out_dup_0[102]), .D (in_int[479]), .C (clk_int)) ;
    FD \reg_out(101)  (.Q (out_dup_0[101]), .D (in_int[480]), .C (clk_int)) ;
    FD \reg_out(100)  (.Q (out_dup_0[100]), .D (in_int[481]), .C (clk_int)) ;
    FD \reg_out(99)  (.Q (out_dup_0[99]), .D (in_int[482]), .C (clk_int)) ;
    FD \reg_out(98)  (.Q (out_dup_0[98]), .D (in_int[483]), .C (clk_int)) ;
    FD \reg_out(97)  (.Q (out_dup_0[97]), .D (in_int[484]), .C (clk_int)) ;
    FD \reg_out(96)  (.Q (out_dup_0[96]), .D (in_int[485]), .C (clk_int)) ;
    FD \reg_out(95)  (.Q (out_dup_0[95]), .D (in_int[486]), .C (clk_int)) ;
    FD \reg_out(94)  (.Q (out_dup_0[94]), .D (in_int[487]), .C (clk_int)) ;
    FD \reg_out(93)  (.Q (out_dup_0[93]), .D (in_int[488]), .C (clk_int)) ;
    FD \reg_out(92)  (.Q (out_dup_0[92]), .D (in_int[489]), .C (clk_int)) ;
    FD \reg_out(91)  (.Q (out_dup_0[91]), .D (in_int[490]), .C (clk_int)) ;
    FD \reg_out(90)  (.Q (out_dup_0[90]), .D (in_int[491]), .C (clk_int)) ;
    FD \reg_out(89)  (.Q (out_dup_0[89]), .D (in_int[492]), .C (clk_int)) ;
    FD \reg_out(88)  (.Q (out_dup_0[88]), .D (in_int[493]), .C (clk_int)) ;
    FD \reg_out(87)  (.Q (out_dup_0[87]), .D (in_int[494]), .C (clk_int)) ;
    FD \reg_out(86)  (.Q (out_dup_0[86]), .D (in_int[495]), .C (clk_int)) ;
    FD \reg_out(85)  (.Q (out_dup_0[85]), .D (in_int[496]), .C (clk_int)) ;
    FD \reg_out(84)  (.Q (out_dup_0[84]), .D (in_int[497]), .C (clk_int)) ;
    FD \reg_out(83)  (.Q (out_dup_0[83]), .D (in_int[498]), .C (clk_int)) ;
    FD \reg_out(82)  (.Q (out_dup_0[82]), .D (in_int[499]), .C (clk_int)) ;
    FD \reg_out(81)  (.Q (out_dup_0[81]), .D (in_int[500]), .C (clk_int)) ;
    FD \reg_out(80)  (.Q (out_dup_0[80]), .D (in_int[501]), .C (clk_int)) ;
    FD \reg_out(79)  (.Q (out_dup_0[79]), .D (in_int[502]), .C (clk_int)) ;
    FD \reg_out(78)  (.Q (out_dup_0[78]), .D (in_int[503]), .C (clk_int)) ;
    FD \reg_out(77)  (.Q (out_dup_0[77]), .D (in_int[504]), .C (clk_int)) ;
    FD \reg_out(76)  (.Q (out_dup_0[76]), .D (in_int[505]), .C (clk_int)) ;
    FD \reg_out(75)  (.Q (out_dup_0[75]), .D (in_int[506]), .C (clk_int)) ;
    FD \reg_out(74)  (.Q (out_dup_0[74]), .D (in_int[507]), .C (clk_int)) ;
    FD \reg_out(73)  (.Q (out_dup_0[73]), .D (in_int[508]), .C (clk_int)) ;
    FD \reg_out(72)  (.Q (out_dup_0[72]), .D (in_int[509]), .C (clk_int)) ;
    FD \reg_out(71)  (.Q (out_dup_0[71]), .D (in_int[510]), .C (clk_int)) ;
    FD \reg_out(70)  (.Q (out_dup_0[70]), .D (in_int[511]), .C (clk_int)) ;
    FD \reg_out(69)  (.Q (out_dup_0[69]), .D (in_int[512]), .C (clk_int)) ;
    FD \reg_out(68)  (.Q (out_dup_0[68]), .D (in_int[513]), .C (clk_int)) ;
    FD \reg_out(67)  (.Q (out_dup_0[67]), .D (in_int[514]), .C (clk_int)) ;
    FD \reg_out(66)  (.Q (out_dup_0[66]), .D (in_int[515]), .C (clk_int)) ;
    FD \reg_out(65)  (.Q (out_dup_0[65]), .D (in_int[516]), .C (clk_int)) ;
    FD \reg_out(64)  (.Q (out_dup_0[64]), .D (in_int[517]), .C (clk_int)) ;
    FD \reg_out(63)  (.Q (out_dup_0[63]), .D (in_int[518]), .C (clk_int)) ;
    FD \reg_out(62)  (.Q (out_dup_0[62]), .D (in_int[519]), .C (clk_int)) ;
    FD \reg_out(61)  (.Q (out_dup_0[61]), .D (in_int[520]), .C (clk_int)) ;
    FD \reg_out(60)  (.Q (out_dup_0[60]), .D (in_int[521]), .C (clk_int)) ;
    FD \reg_out(59)  (.Q (out_dup_0[59]), .D (in_int[522]), .C (clk_int)) ;
    FD \reg_out(58)  (.Q (out_dup_0[58]), .D (in_int[523]), .C (clk_int)) ;
    FD \reg_out(57)  (.Q (out_dup_0[57]), .D (in_int[524]), .C (clk_int)) ;
    FD \reg_out(56)  (.Q (out_dup_0[56]), .D (in_int[525]), .C (clk_int)) ;
    FD \reg_out(55)  (.Q (out_dup_0[55]), .D (in_int[526]), .C (clk_int)) ;
    FD \reg_out(54)  (.Q (out_dup_0[54]), .D (in_int[527]), .C (clk_int)) ;
    FD \reg_out(53)  (.Q (out_dup_0[53]), .D (in_int[528]), .C (clk_int)) ;
    FD \reg_out(52)  (.Q (out_dup_0[52]), .D (in_int[529]), .C (clk_int)) ;
    FD \reg_out(51)  (.Q (out_dup_0[51]), .D (in_int[530]), .C (clk_int)) ;
    FD \reg_out(50)  (.Q (out_dup_0[50]), .D (in_int[531]), .C (clk_int)) ;
    FD \reg_out(49)  (.Q (out_dup_0[49]), .D (in_int[532]), .C (clk_int)) ;
    FD \reg_out(48)  (.Q (out_dup_0[48]), .D (in_int[533]), .C (clk_int)) ;
    FD \reg_out(47)  (.Q (out_dup_0[47]), .D (in_int[534]), .C (clk_int)) ;
    FD \reg_out(46)  (.Q (out_dup_0[46]), .D (in_int[535]), .C (clk_int)) ;
    FD \reg_out(45)  (.Q (out_dup_0[45]), .D (in_int[536]), .C (clk_int)) ;
    FD \reg_out(44)  (.Q (out_dup_0[44]), .D (in_int[537]), .C (clk_int)) ;
    FD \reg_out(43)  (.Q (out_dup_0[43]), .D (in_int[538]), .C (clk_int)) ;
    FD \reg_out(42)  (.Q (out_dup_0[42]), .D (in_int[539]), .C (clk_int)) ;
    FD \reg_out(41)  (.Q (out_dup_0[41]), .D (in_int[540]), .C (clk_int)) ;
    FD \reg_out(40)  (.Q (out_dup_0[40]), .D (in_int[541]), .C (clk_int)) ;
    FD \reg_out(39)  (.Q (out_dup_0[39]), .D (in_int[542]), .C (clk_int)) ;
    FD \reg_out(38)  (.Q (out_dup_0[38]), .D (in_int[543]), .C (clk_int)) ;
    FD \reg_out(37)  (.Q (out_dup_0[37]), .D (in_int[544]), .C (clk_int)) ;
    FD \reg_out(36)  (.Q (out_dup_0[36]), .D (in_int[545]), .C (clk_int)) ;
    FD \reg_out(35)  (.Q (out_dup_0[35]), .D (in_int[546]), .C (clk_int)) ;
    FD \reg_out(34)  (.Q (out_dup_0[34]), .D (in_int[547]), .C (clk_int)) ;
    FD \reg_out(33)  (.Q (out_dup_0[33]), .D (in_int[548]), .C (clk_int)) ;
    FD \reg_out(32)  (.Q (out_dup_0[32]), .D (in_int[549]), .C (clk_int)) ;
    FD \reg_out(31)  (.Q (out_dup_0[31]), .D (in_int[550]), .C (clk_int)) ;
    FD \reg_out(30)  (.Q (out_dup_0[30]), .D (in_int[551]), .C (clk_int)) ;
    FD \reg_out(29)  (.Q (out_dup_0[29]), .D (in_int[552]), .C (clk_int)) ;
    FD \reg_out(28)  (.Q (out_dup_0[28]), .D (in_int[553]), .C (clk_int)) ;
    FD \reg_out(27)  (.Q (out_dup_0[27]), .D (in_int[554]), .C (clk_int)) ;
    FD \reg_out(26)  (.Q (out_dup_0[26]), .D (in_int[555]), .C (clk_int)) ;
    FD \reg_out(25)  (.Q (out_dup_0[25]), .D (in_int[556]), .C (clk_int)) ;
    FD \reg_out(24)  (.Q (out_dup_0[24]), .D (in_int[557]), .C (clk_int)) ;
    FD \reg_out(23)  (.Q (out_dup_0[23]), .D (in_int[558]), .C (clk_int)) ;
    FD \reg_out(22)  (.Q (out_dup_0[22]), .D (in_int[559]), .C (clk_int)) ;
    FD \reg_out(21)  (.Q (out_dup_0[21]), .D (in_int[560]), .C (clk_int)) ;
    FD \reg_out(20)  (.Q (out_dup_0[20]), .D (in_int[561]), .C (clk_int)) ;
    FD \reg_out(19)  (.Q (out_dup_0[19]), .D (in_int[562]), .C (clk_int)) ;
    FD \reg_out(18)  (.Q (out_dup_0[18]), .D (in_int[563]), .C (clk_int)) ;
    FD \reg_out(17)  (.Q (out_dup_0[17]), .D (in_int[564]), .C (clk_int)) ;
    FD \reg_out(16)  (.Q (out_dup_0[16]), .D (in_int[565]), .C (clk_int)) ;
    FD \reg_out(15)  (.Q (out_dup_0[15]), .D (in_int[566]), .C (clk_int)) ;
    FD \reg_out(14)  (.Q (out_dup_0[14]), .D (in_int[567]), .C (clk_int)) ;
    FD \reg_out(13)  (.Q (out_dup_0[13]), .D (in_int[568]), .C (clk_int)) ;
    FD \reg_out(12)  (.Q (out_dup_0[12]), .D (in_int[569]), .C (clk_int)) ;
    FD \reg_out(11)  (.Q (out_dup_0[11]), .D (in_int[570]), .C (clk_int)) ;
    FD \reg_out(10)  (.Q (out_dup_0[10]), .D (in_int[571]), .C (clk_int)) ;
    FD \reg_out(9)  (.Q (out_dup_0[9]), .D (in_int[572]), .C (clk_int)) ;
    FD \reg_out(8)  (.Q (out_dup_0[8]), .D (in_int[573]), .C (clk_int)) ;
    FD \reg_out(7)  (.Q (out_dup_0[7]), .D (in_int[574]), .C (clk_int)) ;
    FD \reg_out(6)  (.Q (out_dup_0[6]), .D (in_int[575]), .C (clk_int)) ;
    FD \reg_out(5)  (.Q (out_dup_0[5]), .D (in_int[576]), .C (clk_int)) ;
    FD \reg_out(4)  (.Q (out_dup_0[4]), .D (in_int[577]), .C (clk_int)) ;
    FD \reg_out(3)  (.Q (out_dup_0[3]), .D (in_int[578]), .C (clk_int)) ;
    FD \reg_out(2)  (.Q (out_dup_0[2]), .D (in_int[579]), .C (clk_int)) ;
    FD \reg_out(1)  (.Q (out_dup_0[1]), .D (in_int[580]), .C (clk_int)) ;
    FD \reg_out(0)  (.Q (out_dup_0[0]), .D (in_int[581]), .C (clk_int)) ;
    BUFGP clk_ibuf (.O (clk_int), .I (clk)) ;
endmodule

