/* memory define and read write by verilog */
/* Reference: https://github.com/jjcarrier/FPGA_2_ShiftReg  */
module memory

endmodule
