// test bench
`timescale 1ns/1ps
module top_tb();
    
    defines_test u0();

endmodule
