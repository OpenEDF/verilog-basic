/**********************************************************************
 * Module definition with ports derived from extern declaration
 *
 * Author: Stuart Sutherland
 *
 * (c) Copyright 2003, Sutherland HDL, Inc. *** ALL RIGHTS RESERVED ***
 * www.sutherland-hdl.com
 *
 * Used with permission in the book, "SystemVerilog for Design"
 *  By Stuart Sutherland, Simon Davidmann, and Peter Flake.
 *  Book copyright: 2003, Kluwer Academic Publishers, Norwell, MA, USA
 *  www.wkap.il, ISBN: 0-4020-7530-8
 *
 * Revision History:
 *   1.00 15 Dec 2003 -- original code, as included in book
 *   1.01 10 Jul 2004 -- cleaned up comments, added expected results
 *                       to output messages
 *
 * Caveat: Expected results displayed for this code example are based
 * on an interpretation of the SystemVerilog 3.1 standard by the code
 * author or authors.  At the time of writing, official SystemVerilog
 * validation suites were not available to validate the example.
 *
 * RIGHT TO USE: This code example, or any portion thereof, may be
 * used and distributed without restriction, provided that this entire
 * comment block is included with the example.
 *
 * DISCLAIMER: THIS CODE EXAMPLE IS PROVIDED "AS IS" WITHOUT WARRANTY
 * OF ANY KIND, EITHER EXPRESS OR IMPLIED, INCLUDING, BUT NOT LIMITED
 * TO WARRANTIES OF MERCHANTABILITY, FITNESS OR CORRECTNESS. IN NO
 * EVENT SHALL THE AUTHOR OR AUTHORS BE LIABLE FOR ANY DAMAGES,
 * INCLUDING INCIDENTAL OR CONSEQUENTIAL DAMAGES, ARISING OUT OF THE
 * USE OF THIS CODE.
 *********************************************************************/


// prototype using Verilog-2001 style
extern module counter #(parameter N = 15)
                        (output logic [N:0] cnt,
                         input  wire  [N:0] d,
                         input  wire        clock,
                                            load
                                            resetN);


module counter ( .* );
  always @(posedge clock, negedge resetN) begin
    if (!resetN)   cnt <= 0;
    else if (load) cnt <= d;
    else           cnt <= cnt + 1;
  end
endmodule

module test;

  logic [3:0] cnt, d;
  bit         clock, load, resetN;

  counter #(.N(3)) dut ( .cnt(cnt),
                         .d(d),
                         .clock(clock),
                         .load(load),
                         .resetN(resetN) );

  initial begin
    $display("\nNo simulation results--just checking that example compiles and elaborates.\n");
    $finish;
  end
endmodule
