//
// Verilog description for cell uni_atm, 
// 02/06/14 03:02:33
//
// Precision RTL Synthesis, 2013a.9//


module uni_atm ( clk, rstN, uni_cell_in, \uni_cell_out_Payload_in(47) , 
                 \uni_cell_out_Payload_in(46) , \uni_cell_out_Payload_in(45) , 
                 \uni_cell_out_Payload_in(44) , \uni_cell_out_Payload_in(43) , 
                 \uni_cell_out_Payload_in(42) , \uni_cell_out_Payload_in(41) , 
                 \uni_cell_out_Payload_in(40) , \uni_cell_out_Payload_in(39) , 
                 \uni_cell_out_Payload_in(38) , \uni_cell_out_Payload_in(37) , 
                 \uni_cell_out_Payload_in(36) , \uni_cell_out_Payload_in(35) , 
                 \uni_cell_out_Payload_in(34) , \uni_cell_out_Payload_in(33) , 
                 \uni_cell_out_Payload_in(32) , \uni_cell_out_Payload_in(31) , 
                 \uni_cell_out_Payload_in(30) , \uni_cell_out_Payload_in(29) , 
                 \uni_cell_out_Payload_in(28) , \uni_cell_out_Payload_in(27) , 
                 \uni_cell_out_Payload_in(26) , \uni_cell_out_Payload_in(25) , 
                 \uni_cell_out_Payload_in(24) , \uni_cell_out_Payload_in(23) , 
                 \uni_cell_out_Payload_in(22) , \uni_cell_out_Payload_in(21) , 
                 \uni_cell_out_Payload_in(20) , \uni_cell_out_Payload_in(19) , 
                 \uni_cell_out_Payload_in(18) , \uni_cell_out_Payload_in(17) , 
                 \uni_cell_out_Payload_in(16) , \uni_cell_out_Payload_in(15) , 
                 \uni_cell_out_Payload_in(14) , \uni_cell_out_Payload_in(13) , 
                 \uni_cell_out_Payload_in(12) , \uni_cell_out_Payload_in(11) , 
                 \uni_cell_out_Payload_in(10) , \uni_cell_out_Payload_in(9) , 
                 \uni_cell_out_Payload_in(8) , \uni_cell_out_Payload_in(7) , 
                 \uni_cell_out_Payload_in(6) , \uni_cell_out_Payload_in(5) , 
                 \uni_cell_out_Payload_in(4) , \uni_cell_out_Payload_in(3) , 
                 \uni_cell_out_Payload_in(2) , \uni_cell_out_Payload_in(1) , 
                 \uni_cell_out_Payload_in(0) , uni_cell_out_HEC_in, 
                 uni_cell_out_CLP_in, uni_cell_out_PTI_in, uni_cell_out_VCI_in, 
                 uni_cell_out_VPI_in, uni_cell_out_GFC_in ) ;

    input clk ;
    input rstN ;
    input [423:0]uni_cell_in ;
    output [7:0]\uni_cell_out_Payload_in(47)  ;
    output [7:0]\uni_cell_out_Payload_in(46)  ;
    output [7:0]\uni_cell_out_Payload_in(45)  ;
    output [7:0]\uni_cell_out_Payload_in(44)  ;
    output [7:0]\uni_cell_out_Payload_in(43)  ;
    output [7:0]\uni_cell_out_Payload_in(42)  ;
    output [7:0]\uni_cell_out_Payload_in(41)  ;
    output [7:0]\uni_cell_out_Payload_in(40)  ;
    output [7:0]\uni_cell_out_Payload_in(39)  ;
    output [7:0]\uni_cell_out_Payload_in(38)  ;
    output [7:0]\uni_cell_out_Payload_in(37)  ;
    output [7:0]\uni_cell_out_Payload_in(36)  ;
    output [7:0]\uni_cell_out_Payload_in(35)  ;
    output [7:0]\uni_cell_out_Payload_in(34)  ;
    output [7:0]\uni_cell_out_Payload_in(33)  ;
    output [7:0]\uni_cell_out_Payload_in(32)  ;
    output [7:0]\uni_cell_out_Payload_in(31)  ;
    output [7:0]\uni_cell_out_Payload_in(30)  ;
    output [7:0]\uni_cell_out_Payload_in(29)  ;
    output [7:0]\uni_cell_out_Payload_in(28)  ;
    output [7:0]\uni_cell_out_Payload_in(27)  ;
    output [7:0]\uni_cell_out_Payload_in(26)  ;
    output [7:0]\uni_cell_out_Payload_in(25)  ;
    output [7:0]\uni_cell_out_Payload_in(24)  ;
    output [7:0]\uni_cell_out_Payload_in(23)  ;
    output [7:0]\uni_cell_out_Payload_in(22)  ;
    output [7:0]\uni_cell_out_Payload_in(21)  ;
    output [7:0]\uni_cell_out_Payload_in(20)  ;
    output [7:0]\uni_cell_out_Payload_in(19)  ;
    output [7:0]\uni_cell_out_Payload_in(18)  ;
    output [7:0]\uni_cell_out_Payload_in(17)  ;
    output [7:0]\uni_cell_out_Payload_in(16)  ;
    output [7:0]\uni_cell_out_Payload_in(15)  ;
    output [7:0]\uni_cell_out_Payload_in(14)  ;
    output [7:0]\uni_cell_out_Payload_in(13)  ;
    output [7:0]\uni_cell_out_Payload_in(12)  ;
    output [7:0]\uni_cell_out_Payload_in(11)  ;
    output [7:0]\uni_cell_out_Payload_in(10)  ;
    output [7:0]\uni_cell_out_Payload_in(9)  ;
    output [7:0]\uni_cell_out_Payload_in(8)  ;
    output [7:0]\uni_cell_out_Payload_in(7)  ;
    output [7:0]\uni_cell_out_Payload_in(6)  ;
    output [7:0]\uni_cell_out_Payload_in(5)  ;
    output [7:0]\uni_cell_out_Payload_in(4)  ;
    output [7:0]\uni_cell_out_Payload_in(3)  ;
    output [7:0]\uni_cell_out_Payload_in(2)  ;
    output [7:0]\uni_cell_out_Payload_in(1)  ;
    output [7:0]\uni_cell_out_Payload_in(0)  ;
    output [7:0]uni_cell_out_HEC_in ;
    output uni_cell_out_CLP_in ;
    output [2:0]uni_cell_out_PTI_in ;
    output [15:0]uni_cell_out_VCI_in ;
    output [7:0]uni_cell_out_VPI_in ;
    output [3:0]uni_cell_out_GFC_in ;

    wire [7:0]uni_cell_out_Payload_in_dup_0;
    wire \uni_cell_out_Payload_in(46)_dup_0(7)  , 
         \uni_cell_out_Payload_in(46)_dup_0(6)  , 
         \uni_cell_out_Payload_in(46)_dup_0(5)  , 
         \uni_cell_out_Payload_in(46)_dup_0(4)  , 
         \uni_cell_out_Payload_in(46)_dup_0(3)  , 
         \uni_cell_out_Payload_in(46)_dup_0(2)  , 
         \uni_cell_out_Payload_in(46)_dup_0(1)  , 
         \uni_cell_out_Payload_in(46)_dup_0(0)  , 
         \uni_cell_out_Payload_in(45)_dup_0(7)  , 
         \uni_cell_out_Payload_in(45)_dup_0(6)  , 
         \uni_cell_out_Payload_in(45)_dup_0(5)  , 
         \uni_cell_out_Payload_in(45)_dup_0(4)  , 
         \uni_cell_out_Payload_in(45)_dup_0(3)  , 
         \uni_cell_out_Payload_in(45)_dup_0(2)  , 
         \uni_cell_out_Payload_in(45)_dup_0(1)  , 
         \uni_cell_out_Payload_in(45)_dup_0(0)  , 
         \uni_cell_out_Payload_in(44)_dup_0(7)  , 
         \uni_cell_out_Payload_in(44)_dup_0(6)  , 
         \uni_cell_out_Payload_in(44)_dup_0(5)  , 
         \uni_cell_out_Payload_in(44)_dup_0(4)  , 
         \uni_cell_out_Payload_in(44)_dup_0(3)  , 
         \uni_cell_out_Payload_in(44)_dup_0(2)  , 
         \uni_cell_out_Payload_in(44)_dup_0(1)  , 
         \uni_cell_out_Payload_in(44)_dup_0(0)  , 
         \uni_cell_out_Payload_in(43)_dup_0(7)  , 
         \uni_cell_out_Payload_in(43)_dup_0(6)  , 
         \uni_cell_out_Payload_in(43)_dup_0(5)  , 
         \uni_cell_out_Payload_in(43)_dup_0(4)  , 
         \uni_cell_out_Payload_in(43)_dup_0(3)  , 
         \uni_cell_out_Payload_in(43)_dup_0(2)  , 
         \uni_cell_out_Payload_in(43)_dup_0(1)  , 
         \uni_cell_out_Payload_in(43)_dup_0(0)  , 
         \uni_cell_out_Payload_in(42)_dup_0(7)  , 
         \uni_cell_out_Payload_in(42)_dup_0(6)  , 
         \uni_cell_out_Payload_in(42)_dup_0(5)  , 
         \uni_cell_out_Payload_in(42)_dup_0(4)  , 
         \uni_cell_out_Payload_in(42)_dup_0(3)  , 
         \uni_cell_out_Payload_in(42)_dup_0(2)  , 
         \uni_cell_out_Payload_in(42)_dup_0(1)  , 
         \uni_cell_out_Payload_in(42)_dup_0(0)  , 
         \uni_cell_out_Payload_in(41)_dup_0(7)  , 
         \uni_cell_out_Payload_in(41)_dup_0(6)  , 
         \uni_cell_out_Payload_in(41)_dup_0(5)  , 
         \uni_cell_out_Payload_in(41)_dup_0(4)  , 
         \uni_cell_out_Payload_in(41)_dup_0(3)  , 
         \uni_cell_out_Payload_in(41)_dup_0(2)  , 
         \uni_cell_out_Payload_in(41)_dup_0(1)  , 
         \uni_cell_out_Payload_in(41)_dup_0(0)  , 
         \uni_cell_out_Payload_in(40)_dup_0(7)  , 
         \uni_cell_out_Payload_in(40)_dup_0(6)  , 
         \uni_cell_out_Payload_in(40)_dup_0(5)  , 
         \uni_cell_out_Payload_in(40)_dup_0(4)  , 
         \uni_cell_out_Payload_in(40)_dup_0(3)  , 
         \uni_cell_out_Payload_in(40)_dup_0(2)  , 
         \uni_cell_out_Payload_in(40)_dup_0(1)  , 
         \uni_cell_out_Payload_in(40)_dup_0(0)  , 
         \uni_cell_out_Payload_in(39)_dup_0(7)  , 
         \uni_cell_out_Payload_in(39)_dup_0(6)  , 
         \uni_cell_out_Payload_in(39)_dup_0(5)  , 
         \uni_cell_out_Payload_in(39)_dup_0(4)  , 
         \uni_cell_out_Payload_in(39)_dup_0(3)  , 
         \uni_cell_out_Payload_in(39)_dup_0(2)  , 
         \uni_cell_out_Payload_in(39)_dup_0(1)  , 
         \uni_cell_out_Payload_in(39)_dup_0(0)  , 
         \uni_cell_out_Payload_in(38)_dup_0(7)  , 
         \uni_cell_out_Payload_in(38)_dup_0(6)  , 
         \uni_cell_out_Payload_in(38)_dup_0(5)  , 
         \uni_cell_out_Payload_in(38)_dup_0(4)  , 
         \uni_cell_out_Payload_in(38)_dup_0(3)  , 
         \uni_cell_out_Payload_in(38)_dup_0(2)  , 
         \uni_cell_out_Payload_in(38)_dup_0(1)  , 
         \uni_cell_out_Payload_in(38)_dup_0(0)  , 
         \uni_cell_out_Payload_in(37)_dup_0(7)  , 
         \uni_cell_out_Payload_in(37)_dup_0(6)  , 
         \uni_cell_out_Payload_in(37)_dup_0(5)  , 
         \uni_cell_out_Payload_in(37)_dup_0(4)  , 
         \uni_cell_out_Payload_in(37)_dup_0(3)  , 
         \uni_cell_out_Payload_in(37)_dup_0(2)  , 
         \uni_cell_out_Payload_in(37)_dup_0(1)  , 
         \uni_cell_out_Payload_in(37)_dup_0(0)  , 
         \uni_cell_out_Payload_in(36)_dup_0(7)  , 
         \uni_cell_out_Payload_in(36)_dup_0(6)  , 
         \uni_cell_out_Payload_in(36)_dup_0(5)  , 
         \uni_cell_out_Payload_in(36)_dup_0(4)  , 
         \uni_cell_out_Payload_in(36)_dup_0(3)  , 
         \uni_cell_out_Payload_in(36)_dup_0(2)  , 
         \uni_cell_out_Payload_in(36)_dup_0(1)  , 
         \uni_cell_out_Payload_in(36)_dup_0(0)  , 
         \uni_cell_out_Payload_in(35)_dup_0(7)  , 
         \uni_cell_out_Payload_in(35)_dup_0(6)  , 
         \uni_cell_out_Payload_in(35)_dup_0(5)  , 
         \uni_cell_out_Payload_in(35)_dup_0(4)  , 
         \uni_cell_out_Payload_in(35)_dup_0(3)  , 
         \uni_cell_out_Payload_in(35)_dup_0(2)  , 
         \uni_cell_out_Payload_in(35)_dup_0(1)  , 
         \uni_cell_out_Payload_in(35)_dup_0(0)  , 
         \uni_cell_out_Payload_in(34)_dup_0(7)  , 
         \uni_cell_out_Payload_in(34)_dup_0(6)  , 
         \uni_cell_out_Payload_in(34)_dup_0(5)  , 
         \uni_cell_out_Payload_in(34)_dup_0(4)  , 
         \uni_cell_out_Payload_in(34)_dup_0(3)  , 
         \uni_cell_out_Payload_in(34)_dup_0(2)  , 
         \uni_cell_out_Payload_in(34)_dup_0(1)  , 
         \uni_cell_out_Payload_in(34)_dup_0(0)  , 
         \uni_cell_out_Payload_in(33)_dup_0(7)  , 
         \uni_cell_out_Payload_in(33)_dup_0(6)  , 
         \uni_cell_out_Payload_in(33)_dup_0(5)  , 
         \uni_cell_out_Payload_in(33)_dup_0(4)  , 
         \uni_cell_out_Payload_in(33)_dup_0(3)  , 
         \uni_cell_out_Payload_in(33)_dup_0(2)  , 
         \uni_cell_out_Payload_in(33)_dup_0(1)  , 
         \uni_cell_out_Payload_in(33)_dup_0(0)  , 
         \uni_cell_out_Payload_in(32)_dup_0(7)  , 
         \uni_cell_out_Payload_in(32)_dup_0(6)  , 
         \uni_cell_out_Payload_in(32)_dup_0(5)  , 
         \uni_cell_out_Payload_in(32)_dup_0(4)  , 
         \uni_cell_out_Payload_in(32)_dup_0(3)  , 
         \uni_cell_out_Payload_in(32)_dup_0(2)  , 
         \uni_cell_out_Payload_in(32)_dup_0(1)  , 
         \uni_cell_out_Payload_in(32)_dup_0(0)  , 
         \uni_cell_out_Payload_in(31)_dup_0(7)  , 
         \uni_cell_out_Payload_in(31)_dup_0(6)  , 
         \uni_cell_out_Payload_in(31)_dup_0(5)  , 
         \uni_cell_out_Payload_in(31)_dup_0(4)  , 
         \uni_cell_out_Payload_in(31)_dup_0(3)  , 
         \uni_cell_out_Payload_in(31)_dup_0(2)  , 
         \uni_cell_out_Payload_in(31)_dup_0(1)  , 
         \uni_cell_out_Payload_in(31)_dup_0(0)  , 
         \uni_cell_out_Payload_in(30)_dup_0(7)  , 
         \uni_cell_out_Payload_in(30)_dup_0(6)  , 
         \uni_cell_out_Payload_in(30)_dup_0(5)  , 
         \uni_cell_out_Payload_in(30)_dup_0(4)  , 
         \uni_cell_out_Payload_in(30)_dup_0(3)  , 
         \uni_cell_out_Payload_in(30)_dup_0(2)  , 
         \uni_cell_out_Payload_in(30)_dup_0(1)  , 
         \uni_cell_out_Payload_in(30)_dup_0(0)  , 
         \uni_cell_out_Payload_in(29)_dup_0(7)  , 
         \uni_cell_out_Payload_in(29)_dup_0(6)  , 
         \uni_cell_out_Payload_in(29)_dup_0(5)  , 
         \uni_cell_out_Payload_in(29)_dup_0(4)  , 
         \uni_cell_out_Payload_in(29)_dup_0(3)  , 
         \uni_cell_out_Payload_in(29)_dup_0(2)  , 
         \uni_cell_out_Payload_in(29)_dup_0(1)  , 
         \uni_cell_out_Payload_in(29)_dup_0(0)  , 
         \uni_cell_out_Payload_in(28)_dup_0(7)  , 
         \uni_cell_out_Payload_in(28)_dup_0(6)  , 
         \uni_cell_out_Payload_in(28)_dup_0(5)  , 
         \uni_cell_out_Payload_in(28)_dup_0(4)  , 
         \uni_cell_out_Payload_in(28)_dup_0(3)  , 
         \uni_cell_out_Payload_in(28)_dup_0(2)  , 
         \uni_cell_out_Payload_in(28)_dup_0(1)  , 
         \uni_cell_out_Payload_in(28)_dup_0(0)  , 
         \uni_cell_out_Payload_in(27)_dup_0(7)  , 
         \uni_cell_out_Payload_in(27)_dup_0(6)  , 
         \uni_cell_out_Payload_in(27)_dup_0(5)  , 
         \uni_cell_out_Payload_in(27)_dup_0(4)  , 
         \uni_cell_out_Payload_in(27)_dup_0(3)  , 
         \uni_cell_out_Payload_in(27)_dup_0(2)  , 
         \uni_cell_out_Payload_in(27)_dup_0(1)  , 
         \uni_cell_out_Payload_in(27)_dup_0(0)  , 
         \uni_cell_out_Payload_in(26)_dup_0(7)  , 
         \uni_cell_out_Payload_in(26)_dup_0(6)  , 
         \uni_cell_out_Payload_in(26)_dup_0(5)  , 
         \uni_cell_out_Payload_in(26)_dup_0(4)  , 
         \uni_cell_out_Payload_in(26)_dup_0(3)  , 
         \uni_cell_out_Payload_in(26)_dup_0(2)  , 
         \uni_cell_out_Payload_in(26)_dup_0(1)  , 
         \uni_cell_out_Payload_in(26)_dup_0(0)  , 
         \uni_cell_out_Payload_in(25)_dup_0(7)  , 
         \uni_cell_out_Payload_in(25)_dup_0(6)  , 
         \uni_cell_out_Payload_in(25)_dup_0(5)  , 
         \uni_cell_out_Payload_in(25)_dup_0(4)  , 
         \uni_cell_out_Payload_in(25)_dup_0(3)  , 
         \uni_cell_out_Payload_in(25)_dup_0(2)  , 
         \uni_cell_out_Payload_in(25)_dup_0(1)  , 
         \uni_cell_out_Payload_in(25)_dup_0(0)  , 
         \uni_cell_out_Payload_in(24)_dup_0(7)  , 
         \uni_cell_out_Payload_in(24)_dup_0(6)  , 
         \uni_cell_out_Payload_in(24)_dup_0(5)  , 
         \uni_cell_out_Payload_in(24)_dup_0(4)  , 
         \uni_cell_out_Payload_in(24)_dup_0(3)  , 
         \uni_cell_out_Payload_in(24)_dup_0(2)  , 
         \uni_cell_out_Payload_in(24)_dup_0(1)  , 
         \uni_cell_out_Payload_in(24)_dup_0(0)  , 
         \uni_cell_out_Payload_in(23)_dup_0(7)  , 
         \uni_cell_out_Payload_in(23)_dup_0(6)  , 
         \uni_cell_out_Payload_in(23)_dup_0(5)  , 
         \uni_cell_out_Payload_in(23)_dup_0(4)  , 
         \uni_cell_out_Payload_in(23)_dup_0(3)  , 
         \uni_cell_out_Payload_in(23)_dup_0(2)  , 
         \uni_cell_out_Payload_in(23)_dup_0(1)  , 
         \uni_cell_out_Payload_in(23)_dup_0(0)  , 
         \uni_cell_out_Payload_in(22)_dup_0(7)  , 
         \uni_cell_out_Payload_in(22)_dup_0(6)  , 
         \uni_cell_out_Payload_in(22)_dup_0(5)  , 
         \uni_cell_out_Payload_in(22)_dup_0(4)  , 
         \uni_cell_out_Payload_in(22)_dup_0(3)  , 
         \uni_cell_out_Payload_in(22)_dup_0(2)  , 
         \uni_cell_out_Payload_in(22)_dup_0(1)  , 
         \uni_cell_out_Payload_in(22)_dup_0(0)  , 
         \uni_cell_out_Payload_in(21)_dup_0(7)  , 
         \uni_cell_out_Payload_in(21)_dup_0(6)  , 
         \uni_cell_out_Payload_in(21)_dup_0(5)  , 
         \uni_cell_out_Payload_in(21)_dup_0(4)  , 
         \uni_cell_out_Payload_in(21)_dup_0(3)  , 
         \uni_cell_out_Payload_in(21)_dup_0(2)  , 
         \uni_cell_out_Payload_in(21)_dup_0(1)  , 
         \uni_cell_out_Payload_in(21)_dup_0(0)  , 
         \uni_cell_out_Payload_in(20)_dup_0(7)  , 
         \uni_cell_out_Payload_in(20)_dup_0(6)  , 
         \uni_cell_out_Payload_in(20)_dup_0(5)  , 
         \uni_cell_out_Payload_in(20)_dup_0(4)  , 
         \uni_cell_out_Payload_in(20)_dup_0(3)  , 
         \uni_cell_out_Payload_in(20)_dup_0(2)  , 
         \uni_cell_out_Payload_in(20)_dup_0(1)  , 
         \uni_cell_out_Payload_in(20)_dup_0(0)  , 
         \uni_cell_out_Payload_in(19)_dup_0(7)  , 
         \uni_cell_out_Payload_in(19)_dup_0(6)  , 
         \uni_cell_out_Payload_in(19)_dup_0(5)  , 
         \uni_cell_out_Payload_in(19)_dup_0(4)  , 
         \uni_cell_out_Payload_in(19)_dup_0(3)  , 
         \uni_cell_out_Payload_in(19)_dup_0(2)  , 
         \uni_cell_out_Payload_in(19)_dup_0(1)  , 
         \uni_cell_out_Payload_in(19)_dup_0(0)  , 
         \uni_cell_out_Payload_in(18)_dup_0(7)  , 
         \uni_cell_out_Payload_in(18)_dup_0(6)  , 
         \uni_cell_out_Payload_in(18)_dup_0(5)  , 
         \uni_cell_out_Payload_in(18)_dup_0(4)  , 
         \uni_cell_out_Payload_in(18)_dup_0(3)  , 
         \uni_cell_out_Payload_in(18)_dup_0(2)  , 
         \uni_cell_out_Payload_in(18)_dup_0(1)  , 
         \uni_cell_out_Payload_in(18)_dup_0(0)  , 
         \uni_cell_out_Payload_in(17)_dup_0(7)  , 
         \uni_cell_out_Payload_in(17)_dup_0(6)  , 
         \uni_cell_out_Payload_in(17)_dup_0(5)  , 
         \uni_cell_out_Payload_in(17)_dup_0(4)  , 
         \uni_cell_out_Payload_in(17)_dup_0(3)  , 
         \uni_cell_out_Payload_in(17)_dup_0(2)  , 
         \uni_cell_out_Payload_in(17)_dup_0(1)  , 
         \uni_cell_out_Payload_in(17)_dup_0(0)  , 
         \uni_cell_out_Payload_in(16)_dup_0(7)  , 
         \uni_cell_out_Payload_in(16)_dup_0(6)  , 
         \uni_cell_out_Payload_in(16)_dup_0(5)  , 
         \uni_cell_out_Payload_in(16)_dup_0(4)  , 
         \uni_cell_out_Payload_in(16)_dup_0(3)  , 
         \uni_cell_out_Payload_in(16)_dup_0(2)  , 
         \uni_cell_out_Payload_in(16)_dup_0(1)  , 
         \uni_cell_out_Payload_in(16)_dup_0(0)  , 
         \uni_cell_out_Payload_in(15)_dup_0(7)  , 
         \uni_cell_out_Payload_in(15)_dup_0(6)  , 
         \uni_cell_out_Payload_in(15)_dup_0(5)  , 
         \uni_cell_out_Payload_in(15)_dup_0(4)  , 
         \uni_cell_out_Payload_in(15)_dup_0(3)  , 
         \uni_cell_out_Payload_in(15)_dup_0(2)  , 
         \uni_cell_out_Payload_in(15)_dup_0(1)  , 
         \uni_cell_out_Payload_in(15)_dup_0(0)  , 
         \uni_cell_out_Payload_in(14)_dup_0(7)  , 
         \uni_cell_out_Payload_in(14)_dup_0(6)  , 
         \uni_cell_out_Payload_in(14)_dup_0(5)  , 
         \uni_cell_out_Payload_in(14)_dup_0(4)  , 
         \uni_cell_out_Payload_in(14)_dup_0(3)  , 
         \uni_cell_out_Payload_in(14)_dup_0(2)  , 
         \uni_cell_out_Payload_in(14)_dup_0(1)  , 
         \uni_cell_out_Payload_in(14)_dup_0(0)  , 
         \uni_cell_out_Payload_in(13)_dup_0(7)  , 
         \uni_cell_out_Payload_in(13)_dup_0(6)  , 
         \uni_cell_out_Payload_in(13)_dup_0(5)  , 
         \uni_cell_out_Payload_in(13)_dup_0(4)  , 
         \uni_cell_out_Payload_in(13)_dup_0(3)  , 
         \uni_cell_out_Payload_in(13)_dup_0(2)  , 
         \uni_cell_out_Payload_in(13)_dup_0(1)  , 
         \uni_cell_out_Payload_in(13)_dup_0(0)  , 
         \uni_cell_out_Payload_in(12)_dup_0(7)  , 
         \uni_cell_out_Payload_in(12)_dup_0(6)  , 
         \uni_cell_out_Payload_in(12)_dup_0(5)  , 
         \uni_cell_out_Payload_in(12)_dup_0(4)  , 
         \uni_cell_out_Payload_in(12)_dup_0(3)  , 
         \uni_cell_out_Payload_in(12)_dup_0(2)  , 
         \uni_cell_out_Payload_in(12)_dup_0(1)  , 
         \uni_cell_out_Payload_in(12)_dup_0(0)  , 
         \uni_cell_out_Payload_in(11)_dup_0(7)  , 
         \uni_cell_out_Payload_in(11)_dup_0(6)  , 
         \uni_cell_out_Payload_in(11)_dup_0(5)  , 
         \uni_cell_out_Payload_in(11)_dup_0(4)  , 
         \uni_cell_out_Payload_in(11)_dup_0(3)  , 
         \uni_cell_out_Payload_in(11)_dup_0(2)  , 
         \uni_cell_out_Payload_in(11)_dup_0(1)  , 
         \uni_cell_out_Payload_in(11)_dup_0(0)  , 
         \uni_cell_out_Payload_in(10)_dup_0(7)  , 
         \uni_cell_out_Payload_in(10)_dup_0(6)  , 
         \uni_cell_out_Payload_in(10)_dup_0(5)  , 
         \uni_cell_out_Payload_in(10)_dup_0(4)  , 
         \uni_cell_out_Payload_in(10)_dup_0(3)  , 
         \uni_cell_out_Payload_in(10)_dup_0(2)  , 
         \uni_cell_out_Payload_in(10)_dup_0(1)  , 
         \uni_cell_out_Payload_in(10)_dup_0(0)  , 
         \uni_cell_out_Payload_in(9)_dup_0(7)  , 
         \uni_cell_out_Payload_in(9)_dup_0(6)  , 
         \uni_cell_out_Payload_in(9)_dup_0(5)  , 
         \uni_cell_out_Payload_in(9)_dup_0(4)  , 
         \uni_cell_out_Payload_in(9)_dup_0(3)  , 
         \uni_cell_out_Payload_in(9)_dup_0(2)  , 
         \uni_cell_out_Payload_in(9)_dup_0(1)  , 
         \uni_cell_out_Payload_in(9)_dup_0(0)  , 
         \uni_cell_out_Payload_in(8)_dup_0(7)  , 
         \uni_cell_out_Payload_in(8)_dup_0(6)  , 
         \uni_cell_out_Payload_in(8)_dup_0(5)  , 
         \uni_cell_out_Payload_in(8)_dup_0(4)  , 
         \uni_cell_out_Payload_in(8)_dup_0(3)  , 
         \uni_cell_out_Payload_in(8)_dup_0(2)  , 
         \uni_cell_out_Payload_in(8)_dup_0(1)  , 
         \uni_cell_out_Payload_in(8)_dup_0(0)  , 
         \uni_cell_out_Payload_in(7)_dup_0(7)  , 
         \uni_cell_out_Payload_in(7)_dup_0(6)  , 
         \uni_cell_out_Payload_in(7)_dup_0(5)  , 
         \uni_cell_out_Payload_in(7)_dup_0(4)  , 
         \uni_cell_out_Payload_in(7)_dup_0(3)  , 
         \uni_cell_out_Payload_in(7)_dup_0(2)  , 
         \uni_cell_out_Payload_in(7)_dup_0(1)  , 
         \uni_cell_out_Payload_in(7)_dup_0(0)  , 
         \uni_cell_out_Payload_in(6)_dup_0(7)  , 
         \uni_cell_out_Payload_in(6)_dup_0(6)  , 
         \uni_cell_out_Payload_in(6)_dup_0(5)  , 
         \uni_cell_out_Payload_in(6)_dup_0(4)  , 
         \uni_cell_out_Payload_in(6)_dup_0(3)  , 
         \uni_cell_out_Payload_in(6)_dup_0(2)  , 
         \uni_cell_out_Payload_in(6)_dup_0(1)  , 
         \uni_cell_out_Payload_in(6)_dup_0(0)  , 
         \uni_cell_out_Payload_in(5)_dup_0(7)  , 
         \uni_cell_out_Payload_in(5)_dup_0(6)  , 
         \uni_cell_out_Payload_in(5)_dup_0(5)  , 
         \uni_cell_out_Payload_in(5)_dup_0(4)  , 
         \uni_cell_out_Payload_in(5)_dup_0(3)  , 
         \uni_cell_out_Payload_in(5)_dup_0(2)  , 
         \uni_cell_out_Payload_in(5)_dup_0(1)  , 
         \uni_cell_out_Payload_in(5)_dup_0(0)  , 
         \uni_cell_out_Payload_in(4)_dup_0(7)  , 
         \uni_cell_out_Payload_in(4)_dup_0(6)  , 
         \uni_cell_out_Payload_in(4)_dup_0(5)  , 
         \uni_cell_out_Payload_in(4)_dup_0(4)  , 
         \uni_cell_out_Payload_in(4)_dup_0(3)  , 
         \uni_cell_out_Payload_in(4)_dup_0(2)  , 
         \uni_cell_out_Payload_in(4)_dup_0(1)  , 
         \uni_cell_out_Payload_in(4)_dup_0(0)  , 
         \uni_cell_out_Payload_in(3)_dup_0(7)  , 
         \uni_cell_out_Payload_in(3)_dup_0(6)  , 
         \uni_cell_out_Payload_in(3)_dup_0(5)  , 
         \uni_cell_out_Payload_in(3)_dup_0(4)  , 
         \uni_cell_out_Payload_in(3)_dup_0(3)  , 
         \uni_cell_out_Payload_in(3)_dup_0(2)  , 
         \uni_cell_out_Payload_in(3)_dup_0(1)  , 
         \uni_cell_out_Payload_in(3)_dup_0(0)  , 
         \uni_cell_out_Payload_in(2)_dup_0(7)  , 
         \uni_cell_out_Payload_in(2)_dup_0(6)  , 
         \uni_cell_out_Payload_in(2)_dup_0(5)  , 
         \uni_cell_out_Payload_in(2)_dup_0(4)  , 
         \uni_cell_out_Payload_in(2)_dup_0(3)  , 
         \uni_cell_out_Payload_in(2)_dup_0(2)  , 
         \uni_cell_out_Payload_in(2)_dup_0(1)  , 
         \uni_cell_out_Payload_in(2)_dup_0(0)  , 
         \uni_cell_out_Payload_in(1)_dup_0(7)  , 
         \uni_cell_out_Payload_in(1)_dup_0(6)  , 
         \uni_cell_out_Payload_in(1)_dup_0(5)  , 
         \uni_cell_out_Payload_in(1)_dup_0(4)  , 
         \uni_cell_out_Payload_in(1)_dup_0(3)  , 
         \uni_cell_out_Payload_in(1)_dup_0(2)  , 
         \uni_cell_out_Payload_in(1)_dup_0(1)  , 
         \uni_cell_out_Payload_in(1)_dup_0(0)  , 
         \uni_cell_out_Payload_in(0)_dup_0(7)  , 
         \uni_cell_out_Payload_in(0)_dup_0(6)  , 
         \uni_cell_out_Payload_in(0)_dup_0(5)  , 
         \uni_cell_out_Payload_in(0)_dup_0(4)  , 
         \uni_cell_out_Payload_in(0)_dup_0(3)  , 
         \uni_cell_out_Payload_in(0)_dup_0(2)  , 
         \uni_cell_out_Payload_in(0)_dup_0(1)  , 
         \uni_cell_out_Payload_in(0)_dup_0(0)  ;
    wire [7:0]uni_cell_out_HEC_in_dup_0;
    wire uni_cell_out_CLP_in_dup_0;
    wire [2:0]uni_cell_out_PTI_in_dup_0;
    wire [15:0]uni_cell_out_VCI_in_dup_0;
    wire [7:0]uni_cell_out_VPI_in_dup_0;
    wire [3:0]uni_cell_out_GFC_in_dup_0;
    wire clk_int, rstN_int;
    wire [423:0]uni_cell_in_int;
    wire not_rstN;



    OBUF \uni_cell_out_GFC_in_obuf(0)  (.O (uni_cell_out_GFC_in[0]), .I (
         uni_cell_out_GFC_in_dup_0[0])) ;
    OBUF \uni_cell_out_GFC_in_obuf(1)  (.O (uni_cell_out_GFC_in[1]), .I (
         uni_cell_out_GFC_in_dup_0[1])) ;
    OBUF \uni_cell_out_GFC_in_obuf(2)  (.O (uni_cell_out_GFC_in[2]), .I (
         uni_cell_out_GFC_in_dup_0[2])) ;
    OBUF \uni_cell_out_GFC_in_obuf(3)  (.O (uni_cell_out_GFC_in[3]), .I (
         uni_cell_out_GFC_in_dup_0[3])) ;
    OBUF \uni_cell_out_VPI_in_obuf(0)  (.O (uni_cell_out_VPI_in[0]), .I (
         uni_cell_out_VPI_in_dup_0[0])) ;
    OBUF \uni_cell_out_VPI_in_obuf(1)  (.O (uni_cell_out_VPI_in[1]), .I (
         uni_cell_out_VPI_in_dup_0[1])) ;
    OBUF \uni_cell_out_VPI_in_obuf(2)  (.O (uni_cell_out_VPI_in[2]), .I (
         uni_cell_out_VPI_in_dup_0[2])) ;
    OBUF \uni_cell_out_VPI_in_obuf(3)  (.O (uni_cell_out_VPI_in[3]), .I (
         uni_cell_out_VPI_in_dup_0[3])) ;
    OBUF \uni_cell_out_VPI_in_obuf(4)  (.O (uni_cell_out_VPI_in[4]), .I (
         uni_cell_out_VPI_in_dup_0[4])) ;
    OBUF \uni_cell_out_VPI_in_obuf(5)  (.O (uni_cell_out_VPI_in[5]), .I (
         uni_cell_out_VPI_in_dup_0[5])) ;
    OBUF \uni_cell_out_VPI_in_obuf(6)  (.O (uni_cell_out_VPI_in[6]), .I (
         uni_cell_out_VPI_in_dup_0[6])) ;
    OBUF \uni_cell_out_VPI_in_obuf(7)  (.O (uni_cell_out_VPI_in[7]), .I (
         uni_cell_out_VPI_in_dup_0[7])) ;
    OBUF \uni_cell_out_VCI_in_obuf(0)  (.O (uni_cell_out_VCI_in[0]), .I (
         uni_cell_out_VCI_in_dup_0[0])) ;
    OBUF \uni_cell_out_VCI_in_obuf(1)  (.O (uni_cell_out_VCI_in[1]), .I (
         uni_cell_out_VCI_in_dup_0[1])) ;
    OBUF \uni_cell_out_VCI_in_obuf(2)  (.O (uni_cell_out_VCI_in[2]), .I (
         uni_cell_out_VCI_in_dup_0[2])) ;
    OBUF \uni_cell_out_VCI_in_obuf(3)  (.O (uni_cell_out_VCI_in[3]), .I (
         uni_cell_out_VCI_in_dup_0[3])) ;
    OBUF \uni_cell_out_VCI_in_obuf(4)  (.O (uni_cell_out_VCI_in[4]), .I (
         uni_cell_out_VCI_in_dup_0[4])) ;
    OBUF \uni_cell_out_VCI_in_obuf(5)  (.O (uni_cell_out_VCI_in[5]), .I (
         uni_cell_out_VCI_in_dup_0[5])) ;
    OBUF \uni_cell_out_VCI_in_obuf(6)  (.O (uni_cell_out_VCI_in[6]), .I (
         uni_cell_out_VCI_in_dup_0[6])) ;
    OBUF \uni_cell_out_VCI_in_obuf(7)  (.O (uni_cell_out_VCI_in[7]), .I (
         uni_cell_out_VCI_in_dup_0[7])) ;
    OBUF \uni_cell_out_VCI_in_obuf(8)  (.O (uni_cell_out_VCI_in[8]), .I (
         uni_cell_out_VCI_in_dup_0[8])) ;
    OBUF \uni_cell_out_VCI_in_obuf(9)  (.O (uni_cell_out_VCI_in[9]), .I (
         uni_cell_out_VCI_in_dup_0[9])) ;
    OBUF \uni_cell_out_VCI_in_obuf(10)  (.O (uni_cell_out_VCI_in[10]), .I (
         uni_cell_out_VCI_in_dup_0[10])) ;
    OBUF \uni_cell_out_VCI_in_obuf(11)  (.O (uni_cell_out_VCI_in[11]), .I (
         uni_cell_out_VCI_in_dup_0[11])) ;
    OBUF \uni_cell_out_VCI_in_obuf(12)  (.O (uni_cell_out_VCI_in[12]), .I (
         uni_cell_out_VCI_in_dup_0[12])) ;
    OBUF \uni_cell_out_VCI_in_obuf(13)  (.O (uni_cell_out_VCI_in[13]), .I (
         uni_cell_out_VCI_in_dup_0[13])) ;
    OBUF \uni_cell_out_VCI_in_obuf(14)  (.O (uni_cell_out_VCI_in[14]), .I (
         uni_cell_out_VCI_in_dup_0[14])) ;
    OBUF \uni_cell_out_VCI_in_obuf(15)  (.O (uni_cell_out_VCI_in[15]), .I (
         uni_cell_out_VCI_in_dup_0[15])) ;
    OBUF \uni_cell_out_PTI_in_obuf(0)  (.O (uni_cell_out_PTI_in[0]), .I (
         uni_cell_out_PTI_in_dup_0[0])) ;
    OBUF \uni_cell_out_PTI_in_obuf(1)  (.O (uni_cell_out_PTI_in[1]), .I (
         uni_cell_out_PTI_in_dup_0[1])) ;
    OBUF \uni_cell_out_PTI_in_obuf(2)  (.O (uni_cell_out_PTI_in[2]), .I (
         uni_cell_out_PTI_in_dup_0[2])) ;
    OBUF uni_cell_out_CLP_in_obuf (.O (uni_cell_out_CLP_in), .I (
         uni_cell_out_CLP_in_dup_0)) ;
    OBUF \uni_cell_out_HEC_in_obuf(0)  (.O (uni_cell_out_HEC_in[0]), .I (
         uni_cell_out_HEC_in_dup_0[0])) ;
    OBUF \uni_cell_out_HEC_in_obuf(1)  (.O (uni_cell_out_HEC_in[1]), .I (
         uni_cell_out_HEC_in_dup_0[1])) ;
    OBUF \uni_cell_out_HEC_in_obuf(2)  (.O (uni_cell_out_HEC_in[2]), .I (
         uni_cell_out_HEC_in_dup_0[2])) ;
    OBUF \uni_cell_out_HEC_in_obuf(3)  (.O (uni_cell_out_HEC_in[3]), .I (
         uni_cell_out_HEC_in_dup_0[3])) ;
    OBUF \uni_cell_out_HEC_in_obuf(4)  (.O (uni_cell_out_HEC_in[4]), .I (
         uni_cell_out_HEC_in_dup_0[4])) ;
    OBUF \uni_cell_out_HEC_in_obuf(5)  (.O (uni_cell_out_HEC_in[5]), .I (
         uni_cell_out_HEC_in_dup_0[5])) ;
    OBUF \uni_cell_out_HEC_in_obuf(6)  (.O (uni_cell_out_HEC_in[6]), .I (
         uni_cell_out_HEC_in_dup_0[6])) ;
    OBUF \uni_cell_out_HEC_in_obuf(7)  (.O (uni_cell_out_HEC_in[7]), .I (
         uni_cell_out_HEC_in_dup_0[7])) ;
    OBUF \uni_cell_out_Payload_in_obuf(0)(0)  (.O (
         \uni_cell_out_Payload_in(0) [0]), .I (
         \uni_cell_out_Payload_in(0)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(0)(1)  (.O (
         \uni_cell_out_Payload_in(0) [1]), .I (
         \uni_cell_out_Payload_in(0)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(0)(2)  (.O (
         \uni_cell_out_Payload_in(0) [2]), .I (
         \uni_cell_out_Payload_in(0)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(0)(3)  (.O (
         \uni_cell_out_Payload_in(0) [3]), .I (
         \uni_cell_out_Payload_in(0)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(0)(4)  (.O (
         \uni_cell_out_Payload_in(0) [4]), .I (
         \uni_cell_out_Payload_in(0)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(0)(5)  (.O (
         \uni_cell_out_Payload_in(0) [5]), .I (
         \uni_cell_out_Payload_in(0)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(0)(6)  (.O (
         \uni_cell_out_Payload_in(0) [6]), .I (
         \uni_cell_out_Payload_in(0)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(0)(7)  (.O (
         \uni_cell_out_Payload_in(0) [7]), .I (
         \uni_cell_out_Payload_in(0)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(1)(0)  (.O (
         \uni_cell_out_Payload_in(1) [0]), .I (
         \uni_cell_out_Payload_in(1)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(1)(1)  (.O (
         \uni_cell_out_Payload_in(1) [1]), .I (
         \uni_cell_out_Payload_in(1)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(1)(2)  (.O (
         \uni_cell_out_Payload_in(1) [2]), .I (
         \uni_cell_out_Payload_in(1)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(1)(3)  (.O (
         \uni_cell_out_Payload_in(1) [3]), .I (
         \uni_cell_out_Payload_in(1)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(1)(4)  (.O (
         \uni_cell_out_Payload_in(1) [4]), .I (
         \uni_cell_out_Payload_in(1)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(1)(5)  (.O (
         \uni_cell_out_Payload_in(1) [5]), .I (
         \uni_cell_out_Payload_in(1)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(1)(6)  (.O (
         \uni_cell_out_Payload_in(1) [6]), .I (
         \uni_cell_out_Payload_in(1)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(1)(7)  (.O (
         \uni_cell_out_Payload_in(1) [7]), .I (
         \uni_cell_out_Payload_in(1)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(2)(0)  (.O (
         \uni_cell_out_Payload_in(2) [0]), .I (
         \uni_cell_out_Payload_in(2)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(2)(1)  (.O (
         \uni_cell_out_Payload_in(2) [1]), .I (
         \uni_cell_out_Payload_in(2)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(2)(2)  (.O (
         \uni_cell_out_Payload_in(2) [2]), .I (
         \uni_cell_out_Payload_in(2)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(2)(3)  (.O (
         \uni_cell_out_Payload_in(2) [3]), .I (
         \uni_cell_out_Payload_in(2)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(2)(4)  (.O (
         \uni_cell_out_Payload_in(2) [4]), .I (
         \uni_cell_out_Payload_in(2)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(2)(5)  (.O (
         \uni_cell_out_Payload_in(2) [5]), .I (
         \uni_cell_out_Payload_in(2)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(2)(6)  (.O (
         \uni_cell_out_Payload_in(2) [6]), .I (
         \uni_cell_out_Payload_in(2)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(2)(7)  (.O (
         \uni_cell_out_Payload_in(2) [7]), .I (
         \uni_cell_out_Payload_in(2)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(3)(0)  (.O (
         \uni_cell_out_Payload_in(3) [0]), .I (
         \uni_cell_out_Payload_in(3)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(3)(1)  (.O (
         \uni_cell_out_Payload_in(3) [1]), .I (
         \uni_cell_out_Payload_in(3)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(3)(2)  (.O (
         \uni_cell_out_Payload_in(3) [2]), .I (
         \uni_cell_out_Payload_in(3)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(3)(3)  (.O (
         \uni_cell_out_Payload_in(3) [3]), .I (
         \uni_cell_out_Payload_in(3)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(3)(4)  (.O (
         \uni_cell_out_Payload_in(3) [4]), .I (
         \uni_cell_out_Payload_in(3)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(3)(5)  (.O (
         \uni_cell_out_Payload_in(3) [5]), .I (
         \uni_cell_out_Payload_in(3)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(3)(6)  (.O (
         \uni_cell_out_Payload_in(3) [6]), .I (
         \uni_cell_out_Payload_in(3)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(3)(7)  (.O (
         \uni_cell_out_Payload_in(3) [7]), .I (
         \uni_cell_out_Payload_in(3)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(4)(0)  (.O (
         \uni_cell_out_Payload_in(4) [0]), .I (
         \uni_cell_out_Payload_in(4)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(4)(1)  (.O (
         \uni_cell_out_Payload_in(4) [1]), .I (
         \uni_cell_out_Payload_in(4)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(4)(2)  (.O (
         \uni_cell_out_Payload_in(4) [2]), .I (
         \uni_cell_out_Payload_in(4)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(4)(3)  (.O (
         \uni_cell_out_Payload_in(4) [3]), .I (
         \uni_cell_out_Payload_in(4)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(4)(4)  (.O (
         \uni_cell_out_Payload_in(4) [4]), .I (
         \uni_cell_out_Payload_in(4)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(4)(5)  (.O (
         \uni_cell_out_Payload_in(4) [5]), .I (
         \uni_cell_out_Payload_in(4)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(4)(6)  (.O (
         \uni_cell_out_Payload_in(4) [6]), .I (
         \uni_cell_out_Payload_in(4)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(4)(7)  (.O (
         \uni_cell_out_Payload_in(4) [7]), .I (
         \uni_cell_out_Payload_in(4)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(5)(0)  (.O (
         \uni_cell_out_Payload_in(5) [0]), .I (
         \uni_cell_out_Payload_in(5)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(5)(1)  (.O (
         \uni_cell_out_Payload_in(5) [1]), .I (
         \uni_cell_out_Payload_in(5)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(5)(2)  (.O (
         \uni_cell_out_Payload_in(5) [2]), .I (
         \uni_cell_out_Payload_in(5)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(5)(3)  (.O (
         \uni_cell_out_Payload_in(5) [3]), .I (
         \uni_cell_out_Payload_in(5)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(5)(4)  (.O (
         \uni_cell_out_Payload_in(5) [4]), .I (
         \uni_cell_out_Payload_in(5)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(5)(5)  (.O (
         \uni_cell_out_Payload_in(5) [5]), .I (
         \uni_cell_out_Payload_in(5)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(5)(6)  (.O (
         \uni_cell_out_Payload_in(5) [6]), .I (
         \uni_cell_out_Payload_in(5)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(5)(7)  (.O (
         \uni_cell_out_Payload_in(5) [7]), .I (
         \uni_cell_out_Payload_in(5)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(6)(0)  (.O (
         \uni_cell_out_Payload_in(6) [0]), .I (
         \uni_cell_out_Payload_in(6)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(6)(1)  (.O (
         \uni_cell_out_Payload_in(6) [1]), .I (
         \uni_cell_out_Payload_in(6)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(6)(2)  (.O (
         \uni_cell_out_Payload_in(6) [2]), .I (
         \uni_cell_out_Payload_in(6)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(6)(3)  (.O (
         \uni_cell_out_Payload_in(6) [3]), .I (
         \uni_cell_out_Payload_in(6)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(6)(4)  (.O (
         \uni_cell_out_Payload_in(6) [4]), .I (
         \uni_cell_out_Payload_in(6)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(6)(5)  (.O (
         \uni_cell_out_Payload_in(6) [5]), .I (
         \uni_cell_out_Payload_in(6)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(6)(6)  (.O (
         \uni_cell_out_Payload_in(6) [6]), .I (
         \uni_cell_out_Payload_in(6)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(6)(7)  (.O (
         \uni_cell_out_Payload_in(6) [7]), .I (
         \uni_cell_out_Payload_in(6)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(7)(0)  (.O (
         \uni_cell_out_Payload_in(7) [0]), .I (
         \uni_cell_out_Payload_in(7)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(7)(1)  (.O (
         \uni_cell_out_Payload_in(7) [1]), .I (
         \uni_cell_out_Payload_in(7)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(7)(2)  (.O (
         \uni_cell_out_Payload_in(7) [2]), .I (
         \uni_cell_out_Payload_in(7)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(7)(3)  (.O (
         \uni_cell_out_Payload_in(7) [3]), .I (
         \uni_cell_out_Payload_in(7)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(7)(4)  (.O (
         \uni_cell_out_Payload_in(7) [4]), .I (
         \uni_cell_out_Payload_in(7)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(7)(5)  (.O (
         \uni_cell_out_Payload_in(7) [5]), .I (
         \uni_cell_out_Payload_in(7)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(7)(6)  (.O (
         \uni_cell_out_Payload_in(7) [6]), .I (
         \uni_cell_out_Payload_in(7)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(7)(7)  (.O (
         \uni_cell_out_Payload_in(7) [7]), .I (
         \uni_cell_out_Payload_in(7)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(8)(0)  (.O (
         \uni_cell_out_Payload_in(8) [0]), .I (
         \uni_cell_out_Payload_in(8)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(8)(1)  (.O (
         \uni_cell_out_Payload_in(8) [1]), .I (
         \uni_cell_out_Payload_in(8)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(8)(2)  (.O (
         \uni_cell_out_Payload_in(8) [2]), .I (
         \uni_cell_out_Payload_in(8)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(8)(3)  (.O (
         \uni_cell_out_Payload_in(8) [3]), .I (
         \uni_cell_out_Payload_in(8)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(8)(4)  (.O (
         \uni_cell_out_Payload_in(8) [4]), .I (
         \uni_cell_out_Payload_in(8)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(8)(5)  (.O (
         \uni_cell_out_Payload_in(8) [5]), .I (
         \uni_cell_out_Payload_in(8)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(8)(6)  (.O (
         \uni_cell_out_Payload_in(8) [6]), .I (
         \uni_cell_out_Payload_in(8)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(8)(7)  (.O (
         \uni_cell_out_Payload_in(8) [7]), .I (
         \uni_cell_out_Payload_in(8)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(9)(0)  (.O (
         \uni_cell_out_Payload_in(9) [0]), .I (
         \uni_cell_out_Payload_in(9)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(9)(1)  (.O (
         \uni_cell_out_Payload_in(9) [1]), .I (
         \uni_cell_out_Payload_in(9)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(9)(2)  (.O (
         \uni_cell_out_Payload_in(9) [2]), .I (
         \uni_cell_out_Payload_in(9)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(9)(3)  (.O (
         \uni_cell_out_Payload_in(9) [3]), .I (
         \uni_cell_out_Payload_in(9)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(9)(4)  (.O (
         \uni_cell_out_Payload_in(9) [4]), .I (
         \uni_cell_out_Payload_in(9)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(9)(5)  (.O (
         \uni_cell_out_Payload_in(9) [5]), .I (
         \uni_cell_out_Payload_in(9)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(9)(6)  (.O (
         \uni_cell_out_Payload_in(9) [6]), .I (
         \uni_cell_out_Payload_in(9)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(9)(7)  (.O (
         \uni_cell_out_Payload_in(9) [7]), .I (
         \uni_cell_out_Payload_in(9)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(10)(0)  (.O (
         \uni_cell_out_Payload_in(10) [0]), .I (
         \uni_cell_out_Payload_in(10)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(10)(1)  (.O (
         \uni_cell_out_Payload_in(10) [1]), .I (
         \uni_cell_out_Payload_in(10)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(10)(2)  (.O (
         \uni_cell_out_Payload_in(10) [2]), .I (
         \uni_cell_out_Payload_in(10)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(10)(3)  (.O (
         \uni_cell_out_Payload_in(10) [3]), .I (
         \uni_cell_out_Payload_in(10)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(10)(4)  (.O (
         \uni_cell_out_Payload_in(10) [4]), .I (
         \uni_cell_out_Payload_in(10)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(10)(5)  (.O (
         \uni_cell_out_Payload_in(10) [5]), .I (
         \uni_cell_out_Payload_in(10)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(10)(6)  (.O (
         \uni_cell_out_Payload_in(10) [6]), .I (
         \uni_cell_out_Payload_in(10)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(10)(7)  (.O (
         \uni_cell_out_Payload_in(10) [7]), .I (
         \uni_cell_out_Payload_in(10)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(11)(0)  (.O (
         \uni_cell_out_Payload_in(11) [0]), .I (
         \uni_cell_out_Payload_in(11)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(11)(1)  (.O (
         \uni_cell_out_Payload_in(11) [1]), .I (
         \uni_cell_out_Payload_in(11)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(11)(2)  (.O (
         \uni_cell_out_Payload_in(11) [2]), .I (
         \uni_cell_out_Payload_in(11)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(11)(3)  (.O (
         \uni_cell_out_Payload_in(11) [3]), .I (
         \uni_cell_out_Payload_in(11)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(11)(4)  (.O (
         \uni_cell_out_Payload_in(11) [4]), .I (
         \uni_cell_out_Payload_in(11)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(11)(5)  (.O (
         \uni_cell_out_Payload_in(11) [5]), .I (
         \uni_cell_out_Payload_in(11)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(11)(6)  (.O (
         \uni_cell_out_Payload_in(11) [6]), .I (
         \uni_cell_out_Payload_in(11)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(11)(7)  (.O (
         \uni_cell_out_Payload_in(11) [7]), .I (
         \uni_cell_out_Payload_in(11)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(12)(0)  (.O (
         \uni_cell_out_Payload_in(12) [0]), .I (
         \uni_cell_out_Payload_in(12)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(12)(1)  (.O (
         \uni_cell_out_Payload_in(12) [1]), .I (
         \uni_cell_out_Payload_in(12)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(12)(2)  (.O (
         \uni_cell_out_Payload_in(12) [2]), .I (
         \uni_cell_out_Payload_in(12)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(12)(3)  (.O (
         \uni_cell_out_Payload_in(12) [3]), .I (
         \uni_cell_out_Payload_in(12)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(12)(4)  (.O (
         \uni_cell_out_Payload_in(12) [4]), .I (
         \uni_cell_out_Payload_in(12)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(12)(5)  (.O (
         \uni_cell_out_Payload_in(12) [5]), .I (
         \uni_cell_out_Payload_in(12)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(12)(6)  (.O (
         \uni_cell_out_Payload_in(12) [6]), .I (
         \uni_cell_out_Payload_in(12)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(12)(7)  (.O (
         \uni_cell_out_Payload_in(12) [7]), .I (
         \uni_cell_out_Payload_in(12)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(13)(0)  (.O (
         \uni_cell_out_Payload_in(13) [0]), .I (
         \uni_cell_out_Payload_in(13)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(13)(1)  (.O (
         \uni_cell_out_Payload_in(13) [1]), .I (
         \uni_cell_out_Payload_in(13)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(13)(2)  (.O (
         \uni_cell_out_Payload_in(13) [2]), .I (
         \uni_cell_out_Payload_in(13)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(13)(3)  (.O (
         \uni_cell_out_Payload_in(13) [3]), .I (
         \uni_cell_out_Payload_in(13)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(13)(4)  (.O (
         \uni_cell_out_Payload_in(13) [4]), .I (
         \uni_cell_out_Payload_in(13)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(13)(5)  (.O (
         \uni_cell_out_Payload_in(13) [5]), .I (
         \uni_cell_out_Payload_in(13)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(13)(6)  (.O (
         \uni_cell_out_Payload_in(13) [6]), .I (
         \uni_cell_out_Payload_in(13)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(13)(7)  (.O (
         \uni_cell_out_Payload_in(13) [7]), .I (
         \uni_cell_out_Payload_in(13)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(14)(0)  (.O (
         \uni_cell_out_Payload_in(14) [0]), .I (
         \uni_cell_out_Payload_in(14)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(14)(1)  (.O (
         \uni_cell_out_Payload_in(14) [1]), .I (
         \uni_cell_out_Payload_in(14)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(14)(2)  (.O (
         \uni_cell_out_Payload_in(14) [2]), .I (
         \uni_cell_out_Payload_in(14)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(14)(3)  (.O (
         \uni_cell_out_Payload_in(14) [3]), .I (
         \uni_cell_out_Payload_in(14)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(14)(4)  (.O (
         \uni_cell_out_Payload_in(14) [4]), .I (
         \uni_cell_out_Payload_in(14)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(14)(5)  (.O (
         \uni_cell_out_Payload_in(14) [5]), .I (
         \uni_cell_out_Payload_in(14)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(14)(6)  (.O (
         \uni_cell_out_Payload_in(14) [6]), .I (
         \uni_cell_out_Payload_in(14)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(14)(7)  (.O (
         \uni_cell_out_Payload_in(14) [7]), .I (
         \uni_cell_out_Payload_in(14)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(15)(0)  (.O (
         \uni_cell_out_Payload_in(15) [0]), .I (
         \uni_cell_out_Payload_in(15)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(15)(1)  (.O (
         \uni_cell_out_Payload_in(15) [1]), .I (
         \uni_cell_out_Payload_in(15)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(15)(2)  (.O (
         \uni_cell_out_Payload_in(15) [2]), .I (
         \uni_cell_out_Payload_in(15)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(15)(3)  (.O (
         \uni_cell_out_Payload_in(15) [3]), .I (
         \uni_cell_out_Payload_in(15)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(15)(4)  (.O (
         \uni_cell_out_Payload_in(15) [4]), .I (
         \uni_cell_out_Payload_in(15)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(15)(5)  (.O (
         \uni_cell_out_Payload_in(15) [5]), .I (
         \uni_cell_out_Payload_in(15)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(15)(6)  (.O (
         \uni_cell_out_Payload_in(15) [6]), .I (
         \uni_cell_out_Payload_in(15)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(15)(7)  (.O (
         \uni_cell_out_Payload_in(15) [7]), .I (
         \uni_cell_out_Payload_in(15)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(16)(0)  (.O (
         \uni_cell_out_Payload_in(16) [0]), .I (
         \uni_cell_out_Payload_in(16)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(16)(1)  (.O (
         \uni_cell_out_Payload_in(16) [1]), .I (
         \uni_cell_out_Payload_in(16)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(16)(2)  (.O (
         \uni_cell_out_Payload_in(16) [2]), .I (
         \uni_cell_out_Payload_in(16)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(16)(3)  (.O (
         \uni_cell_out_Payload_in(16) [3]), .I (
         \uni_cell_out_Payload_in(16)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(16)(4)  (.O (
         \uni_cell_out_Payload_in(16) [4]), .I (
         \uni_cell_out_Payload_in(16)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(16)(5)  (.O (
         \uni_cell_out_Payload_in(16) [5]), .I (
         \uni_cell_out_Payload_in(16)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(16)(6)  (.O (
         \uni_cell_out_Payload_in(16) [6]), .I (
         \uni_cell_out_Payload_in(16)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(16)(7)  (.O (
         \uni_cell_out_Payload_in(16) [7]), .I (
         \uni_cell_out_Payload_in(16)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(17)(0)  (.O (
         \uni_cell_out_Payload_in(17) [0]), .I (
         \uni_cell_out_Payload_in(17)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(17)(1)  (.O (
         \uni_cell_out_Payload_in(17) [1]), .I (
         \uni_cell_out_Payload_in(17)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(17)(2)  (.O (
         \uni_cell_out_Payload_in(17) [2]), .I (
         \uni_cell_out_Payload_in(17)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(17)(3)  (.O (
         \uni_cell_out_Payload_in(17) [3]), .I (
         \uni_cell_out_Payload_in(17)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(17)(4)  (.O (
         \uni_cell_out_Payload_in(17) [4]), .I (
         \uni_cell_out_Payload_in(17)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(17)(5)  (.O (
         \uni_cell_out_Payload_in(17) [5]), .I (
         \uni_cell_out_Payload_in(17)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(17)(6)  (.O (
         \uni_cell_out_Payload_in(17) [6]), .I (
         \uni_cell_out_Payload_in(17)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(17)(7)  (.O (
         \uni_cell_out_Payload_in(17) [7]), .I (
         \uni_cell_out_Payload_in(17)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(18)(0)  (.O (
         \uni_cell_out_Payload_in(18) [0]), .I (
         \uni_cell_out_Payload_in(18)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(18)(1)  (.O (
         \uni_cell_out_Payload_in(18) [1]), .I (
         \uni_cell_out_Payload_in(18)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(18)(2)  (.O (
         \uni_cell_out_Payload_in(18) [2]), .I (
         \uni_cell_out_Payload_in(18)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(18)(3)  (.O (
         \uni_cell_out_Payload_in(18) [3]), .I (
         \uni_cell_out_Payload_in(18)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(18)(4)  (.O (
         \uni_cell_out_Payload_in(18) [4]), .I (
         \uni_cell_out_Payload_in(18)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(18)(5)  (.O (
         \uni_cell_out_Payload_in(18) [5]), .I (
         \uni_cell_out_Payload_in(18)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(18)(6)  (.O (
         \uni_cell_out_Payload_in(18) [6]), .I (
         \uni_cell_out_Payload_in(18)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(18)(7)  (.O (
         \uni_cell_out_Payload_in(18) [7]), .I (
         \uni_cell_out_Payload_in(18)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(19)(0)  (.O (
         \uni_cell_out_Payload_in(19) [0]), .I (
         \uni_cell_out_Payload_in(19)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(19)(1)  (.O (
         \uni_cell_out_Payload_in(19) [1]), .I (
         \uni_cell_out_Payload_in(19)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(19)(2)  (.O (
         \uni_cell_out_Payload_in(19) [2]), .I (
         \uni_cell_out_Payload_in(19)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(19)(3)  (.O (
         \uni_cell_out_Payload_in(19) [3]), .I (
         \uni_cell_out_Payload_in(19)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(19)(4)  (.O (
         \uni_cell_out_Payload_in(19) [4]), .I (
         \uni_cell_out_Payload_in(19)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(19)(5)  (.O (
         \uni_cell_out_Payload_in(19) [5]), .I (
         \uni_cell_out_Payload_in(19)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(19)(6)  (.O (
         \uni_cell_out_Payload_in(19) [6]), .I (
         \uni_cell_out_Payload_in(19)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(19)(7)  (.O (
         \uni_cell_out_Payload_in(19) [7]), .I (
         \uni_cell_out_Payload_in(19)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(20)(0)  (.O (
         \uni_cell_out_Payload_in(20) [0]), .I (
         \uni_cell_out_Payload_in(20)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(20)(1)  (.O (
         \uni_cell_out_Payload_in(20) [1]), .I (
         \uni_cell_out_Payload_in(20)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(20)(2)  (.O (
         \uni_cell_out_Payload_in(20) [2]), .I (
         \uni_cell_out_Payload_in(20)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(20)(3)  (.O (
         \uni_cell_out_Payload_in(20) [3]), .I (
         \uni_cell_out_Payload_in(20)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(20)(4)  (.O (
         \uni_cell_out_Payload_in(20) [4]), .I (
         \uni_cell_out_Payload_in(20)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(20)(5)  (.O (
         \uni_cell_out_Payload_in(20) [5]), .I (
         \uni_cell_out_Payload_in(20)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(20)(6)  (.O (
         \uni_cell_out_Payload_in(20) [6]), .I (
         \uni_cell_out_Payload_in(20)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(20)(7)  (.O (
         \uni_cell_out_Payload_in(20) [7]), .I (
         \uni_cell_out_Payload_in(20)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(21)(0)  (.O (
         \uni_cell_out_Payload_in(21) [0]), .I (
         \uni_cell_out_Payload_in(21)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(21)(1)  (.O (
         \uni_cell_out_Payload_in(21) [1]), .I (
         \uni_cell_out_Payload_in(21)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(21)(2)  (.O (
         \uni_cell_out_Payload_in(21) [2]), .I (
         \uni_cell_out_Payload_in(21)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(21)(3)  (.O (
         \uni_cell_out_Payload_in(21) [3]), .I (
         \uni_cell_out_Payload_in(21)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(21)(4)  (.O (
         \uni_cell_out_Payload_in(21) [4]), .I (
         \uni_cell_out_Payload_in(21)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(21)(5)  (.O (
         \uni_cell_out_Payload_in(21) [5]), .I (
         \uni_cell_out_Payload_in(21)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(21)(6)  (.O (
         \uni_cell_out_Payload_in(21) [6]), .I (
         \uni_cell_out_Payload_in(21)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(21)(7)  (.O (
         \uni_cell_out_Payload_in(21) [7]), .I (
         \uni_cell_out_Payload_in(21)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(22)(0)  (.O (
         \uni_cell_out_Payload_in(22) [0]), .I (
         \uni_cell_out_Payload_in(22)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(22)(1)  (.O (
         \uni_cell_out_Payload_in(22) [1]), .I (
         \uni_cell_out_Payload_in(22)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(22)(2)  (.O (
         \uni_cell_out_Payload_in(22) [2]), .I (
         \uni_cell_out_Payload_in(22)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(22)(3)  (.O (
         \uni_cell_out_Payload_in(22) [3]), .I (
         \uni_cell_out_Payload_in(22)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(22)(4)  (.O (
         \uni_cell_out_Payload_in(22) [4]), .I (
         \uni_cell_out_Payload_in(22)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(22)(5)  (.O (
         \uni_cell_out_Payload_in(22) [5]), .I (
         \uni_cell_out_Payload_in(22)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(22)(6)  (.O (
         \uni_cell_out_Payload_in(22) [6]), .I (
         \uni_cell_out_Payload_in(22)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(22)(7)  (.O (
         \uni_cell_out_Payload_in(22) [7]), .I (
         \uni_cell_out_Payload_in(22)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(23)(0)  (.O (
         \uni_cell_out_Payload_in(23) [0]), .I (
         \uni_cell_out_Payload_in(23)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(23)(1)  (.O (
         \uni_cell_out_Payload_in(23) [1]), .I (
         \uni_cell_out_Payload_in(23)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(23)(2)  (.O (
         \uni_cell_out_Payload_in(23) [2]), .I (
         \uni_cell_out_Payload_in(23)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(23)(3)  (.O (
         \uni_cell_out_Payload_in(23) [3]), .I (
         \uni_cell_out_Payload_in(23)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(23)(4)  (.O (
         \uni_cell_out_Payload_in(23) [4]), .I (
         \uni_cell_out_Payload_in(23)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(23)(5)  (.O (
         \uni_cell_out_Payload_in(23) [5]), .I (
         \uni_cell_out_Payload_in(23)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(23)(6)  (.O (
         \uni_cell_out_Payload_in(23) [6]), .I (
         \uni_cell_out_Payload_in(23)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(23)(7)  (.O (
         \uni_cell_out_Payload_in(23) [7]), .I (
         \uni_cell_out_Payload_in(23)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(24)(0)  (.O (
         \uni_cell_out_Payload_in(24) [0]), .I (
         \uni_cell_out_Payload_in(24)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(24)(1)  (.O (
         \uni_cell_out_Payload_in(24) [1]), .I (
         \uni_cell_out_Payload_in(24)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(24)(2)  (.O (
         \uni_cell_out_Payload_in(24) [2]), .I (
         \uni_cell_out_Payload_in(24)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(24)(3)  (.O (
         \uni_cell_out_Payload_in(24) [3]), .I (
         \uni_cell_out_Payload_in(24)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(24)(4)  (.O (
         \uni_cell_out_Payload_in(24) [4]), .I (
         \uni_cell_out_Payload_in(24)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(24)(5)  (.O (
         \uni_cell_out_Payload_in(24) [5]), .I (
         \uni_cell_out_Payload_in(24)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(24)(6)  (.O (
         \uni_cell_out_Payload_in(24) [6]), .I (
         \uni_cell_out_Payload_in(24)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(24)(7)  (.O (
         \uni_cell_out_Payload_in(24) [7]), .I (
         \uni_cell_out_Payload_in(24)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(25)(0)  (.O (
         \uni_cell_out_Payload_in(25) [0]), .I (
         \uni_cell_out_Payload_in(25)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(25)(1)  (.O (
         \uni_cell_out_Payload_in(25) [1]), .I (
         \uni_cell_out_Payload_in(25)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(25)(2)  (.O (
         \uni_cell_out_Payload_in(25) [2]), .I (
         \uni_cell_out_Payload_in(25)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(25)(3)  (.O (
         \uni_cell_out_Payload_in(25) [3]), .I (
         \uni_cell_out_Payload_in(25)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(25)(4)  (.O (
         \uni_cell_out_Payload_in(25) [4]), .I (
         \uni_cell_out_Payload_in(25)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(25)(5)  (.O (
         \uni_cell_out_Payload_in(25) [5]), .I (
         \uni_cell_out_Payload_in(25)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(25)(6)  (.O (
         \uni_cell_out_Payload_in(25) [6]), .I (
         \uni_cell_out_Payload_in(25)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(25)(7)  (.O (
         \uni_cell_out_Payload_in(25) [7]), .I (
         \uni_cell_out_Payload_in(25)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(26)(0)  (.O (
         \uni_cell_out_Payload_in(26) [0]), .I (
         \uni_cell_out_Payload_in(26)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(26)(1)  (.O (
         \uni_cell_out_Payload_in(26) [1]), .I (
         \uni_cell_out_Payload_in(26)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(26)(2)  (.O (
         \uni_cell_out_Payload_in(26) [2]), .I (
         \uni_cell_out_Payload_in(26)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(26)(3)  (.O (
         \uni_cell_out_Payload_in(26) [3]), .I (
         \uni_cell_out_Payload_in(26)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(26)(4)  (.O (
         \uni_cell_out_Payload_in(26) [4]), .I (
         \uni_cell_out_Payload_in(26)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(26)(5)  (.O (
         \uni_cell_out_Payload_in(26) [5]), .I (
         \uni_cell_out_Payload_in(26)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(26)(6)  (.O (
         \uni_cell_out_Payload_in(26) [6]), .I (
         \uni_cell_out_Payload_in(26)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(26)(7)  (.O (
         \uni_cell_out_Payload_in(26) [7]), .I (
         \uni_cell_out_Payload_in(26)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(27)(0)  (.O (
         \uni_cell_out_Payload_in(27) [0]), .I (
         \uni_cell_out_Payload_in(27)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(27)(1)  (.O (
         \uni_cell_out_Payload_in(27) [1]), .I (
         \uni_cell_out_Payload_in(27)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(27)(2)  (.O (
         \uni_cell_out_Payload_in(27) [2]), .I (
         \uni_cell_out_Payload_in(27)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(27)(3)  (.O (
         \uni_cell_out_Payload_in(27) [3]), .I (
         \uni_cell_out_Payload_in(27)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(27)(4)  (.O (
         \uni_cell_out_Payload_in(27) [4]), .I (
         \uni_cell_out_Payload_in(27)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(27)(5)  (.O (
         \uni_cell_out_Payload_in(27) [5]), .I (
         \uni_cell_out_Payload_in(27)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(27)(6)  (.O (
         \uni_cell_out_Payload_in(27) [6]), .I (
         \uni_cell_out_Payload_in(27)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(27)(7)  (.O (
         \uni_cell_out_Payload_in(27) [7]), .I (
         \uni_cell_out_Payload_in(27)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(28)(0)  (.O (
         \uni_cell_out_Payload_in(28) [0]), .I (
         \uni_cell_out_Payload_in(28)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(28)(1)  (.O (
         \uni_cell_out_Payload_in(28) [1]), .I (
         \uni_cell_out_Payload_in(28)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(28)(2)  (.O (
         \uni_cell_out_Payload_in(28) [2]), .I (
         \uni_cell_out_Payload_in(28)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(28)(3)  (.O (
         \uni_cell_out_Payload_in(28) [3]), .I (
         \uni_cell_out_Payload_in(28)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(28)(4)  (.O (
         \uni_cell_out_Payload_in(28) [4]), .I (
         \uni_cell_out_Payload_in(28)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(28)(5)  (.O (
         \uni_cell_out_Payload_in(28) [5]), .I (
         \uni_cell_out_Payload_in(28)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(28)(6)  (.O (
         \uni_cell_out_Payload_in(28) [6]), .I (
         \uni_cell_out_Payload_in(28)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(28)(7)  (.O (
         \uni_cell_out_Payload_in(28) [7]), .I (
         \uni_cell_out_Payload_in(28)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(29)(0)  (.O (
         \uni_cell_out_Payload_in(29) [0]), .I (
         \uni_cell_out_Payload_in(29)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(29)(1)  (.O (
         \uni_cell_out_Payload_in(29) [1]), .I (
         \uni_cell_out_Payload_in(29)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(29)(2)  (.O (
         \uni_cell_out_Payload_in(29) [2]), .I (
         \uni_cell_out_Payload_in(29)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(29)(3)  (.O (
         \uni_cell_out_Payload_in(29) [3]), .I (
         \uni_cell_out_Payload_in(29)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(29)(4)  (.O (
         \uni_cell_out_Payload_in(29) [4]), .I (
         \uni_cell_out_Payload_in(29)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(29)(5)  (.O (
         \uni_cell_out_Payload_in(29) [5]), .I (
         \uni_cell_out_Payload_in(29)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(29)(6)  (.O (
         \uni_cell_out_Payload_in(29) [6]), .I (
         \uni_cell_out_Payload_in(29)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(29)(7)  (.O (
         \uni_cell_out_Payload_in(29) [7]), .I (
         \uni_cell_out_Payload_in(29)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(30)(0)  (.O (
         \uni_cell_out_Payload_in(30) [0]), .I (
         \uni_cell_out_Payload_in(30)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(30)(1)  (.O (
         \uni_cell_out_Payload_in(30) [1]), .I (
         \uni_cell_out_Payload_in(30)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(30)(2)  (.O (
         \uni_cell_out_Payload_in(30) [2]), .I (
         \uni_cell_out_Payload_in(30)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(30)(3)  (.O (
         \uni_cell_out_Payload_in(30) [3]), .I (
         \uni_cell_out_Payload_in(30)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(30)(4)  (.O (
         \uni_cell_out_Payload_in(30) [4]), .I (
         \uni_cell_out_Payload_in(30)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(30)(5)  (.O (
         \uni_cell_out_Payload_in(30) [5]), .I (
         \uni_cell_out_Payload_in(30)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(30)(6)  (.O (
         \uni_cell_out_Payload_in(30) [6]), .I (
         \uni_cell_out_Payload_in(30)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(30)(7)  (.O (
         \uni_cell_out_Payload_in(30) [7]), .I (
         \uni_cell_out_Payload_in(30)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(31)(0)  (.O (
         \uni_cell_out_Payload_in(31) [0]), .I (
         \uni_cell_out_Payload_in(31)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(31)(1)  (.O (
         \uni_cell_out_Payload_in(31) [1]), .I (
         \uni_cell_out_Payload_in(31)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(31)(2)  (.O (
         \uni_cell_out_Payload_in(31) [2]), .I (
         \uni_cell_out_Payload_in(31)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(31)(3)  (.O (
         \uni_cell_out_Payload_in(31) [3]), .I (
         \uni_cell_out_Payload_in(31)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(31)(4)  (.O (
         \uni_cell_out_Payload_in(31) [4]), .I (
         \uni_cell_out_Payload_in(31)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(31)(5)  (.O (
         \uni_cell_out_Payload_in(31) [5]), .I (
         \uni_cell_out_Payload_in(31)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(31)(6)  (.O (
         \uni_cell_out_Payload_in(31) [6]), .I (
         \uni_cell_out_Payload_in(31)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(31)(7)  (.O (
         \uni_cell_out_Payload_in(31) [7]), .I (
         \uni_cell_out_Payload_in(31)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(32)(0)  (.O (
         \uni_cell_out_Payload_in(32) [0]), .I (
         \uni_cell_out_Payload_in(32)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(32)(1)  (.O (
         \uni_cell_out_Payload_in(32) [1]), .I (
         \uni_cell_out_Payload_in(32)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(32)(2)  (.O (
         \uni_cell_out_Payload_in(32) [2]), .I (
         \uni_cell_out_Payload_in(32)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(32)(3)  (.O (
         \uni_cell_out_Payload_in(32) [3]), .I (
         \uni_cell_out_Payload_in(32)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(32)(4)  (.O (
         \uni_cell_out_Payload_in(32) [4]), .I (
         \uni_cell_out_Payload_in(32)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(32)(5)  (.O (
         \uni_cell_out_Payload_in(32) [5]), .I (
         \uni_cell_out_Payload_in(32)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(32)(6)  (.O (
         \uni_cell_out_Payload_in(32) [6]), .I (
         \uni_cell_out_Payload_in(32)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(32)(7)  (.O (
         \uni_cell_out_Payload_in(32) [7]), .I (
         \uni_cell_out_Payload_in(32)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(33)(0)  (.O (
         \uni_cell_out_Payload_in(33) [0]), .I (
         \uni_cell_out_Payload_in(33)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(33)(1)  (.O (
         \uni_cell_out_Payload_in(33) [1]), .I (
         \uni_cell_out_Payload_in(33)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(33)(2)  (.O (
         \uni_cell_out_Payload_in(33) [2]), .I (
         \uni_cell_out_Payload_in(33)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(33)(3)  (.O (
         \uni_cell_out_Payload_in(33) [3]), .I (
         \uni_cell_out_Payload_in(33)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(33)(4)  (.O (
         \uni_cell_out_Payload_in(33) [4]), .I (
         \uni_cell_out_Payload_in(33)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(33)(5)  (.O (
         \uni_cell_out_Payload_in(33) [5]), .I (
         \uni_cell_out_Payload_in(33)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(33)(6)  (.O (
         \uni_cell_out_Payload_in(33) [6]), .I (
         \uni_cell_out_Payload_in(33)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(33)(7)  (.O (
         \uni_cell_out_Payload_in(33) [7]), .I (
         \uni_cell_out_Payload_in(33)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(34)(0)  (.O (
         \uni_cell_out_Payload_in(34) [0]), .I (
         \uni_cell_out_Payload_in(34)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(34)(1)  (.O (
         \uni_cell_out_Payload_in(34) [1]), .I (
         \uni_cell_out_Payload_in(34)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(34)(2)  (.O (
         \uni_cell_out_Payload_in(34) [2]), .I (
         \uni_cell_out_Payload_in(34)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(34)(3)  (.O (
         \uni_cell_out_Payload_in(34) [3]), .I (
         \uni_cell_out_Payload_in(34)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(34)(4)  (.O (
         \uni_cell_out_Payload_in(34) [4]), .I (
         \uni_cell_out_Payload_in(34)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(34)(5)  (.O (
         \uni_cell_out_Payload_in(34) [5]), .I (
         \uni_cell_out_Payload_in(34)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(34)(6)  (.O (
         \uni_cell_out_Payload_in(34) [6]), .I (
         \uni_cell_out_Payload_in(34)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(34)(7)  (.O (
         \uni_cell_out_Payload_in(34) [7]), .I (
         \uni_cell_out_Payload_in(34)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(35)(0)  (.O (
         \uni_cell_out_Payload_in(35) [0]), .I (
         \uni_cell_out_Payload_in(35)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(35)(1)  (.O (
         \uni_cell_out_Payload_in(35) [1]), .I (
         \uni_cell_out_Payload_in(35)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(35)(2)  (.O (
         \uni_cell_out_Payload_in(35) [2]), .I (
         \uni_cell_out_Payload_in(35)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(35)(3)  (.O (
         \uni_cell_out_Payload_in(35) [3]), .I (
         \uni_cell_out_Payload_in(35)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(35)(4)  (.O (
         \uni_cell_out_Payload_in(35) [4]), .I (
         \uni_cell_out_Payload_in(35)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(35)(5)  (.O (
         \uni_cell_out_Payload_in(35) [5]), .I (
         \uni_cell_out_Payload_in(35)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(35)(6)  (.O (
         \uni_cell_out_Payload_in(35) [6]), .I (
         \uni_cell_out_Payload_in(35)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(35)(7)  (.O (
         \uni_cell_out_Payload_in(35) [7]), .I (
         \uni_cell_out_Payload_in(35)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(36)(0)  (.O (
         \uni_cell_out_Payload_in(36) [0]), .I (
         \uni_cell_out_Payload_in(36)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(36)(1)  (.O (
         \uni_cell_out_Payload_in(36) [1]), .I (
         \uni_cell_out_Payload_in(36)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(36)(2)  (.O (
         \uni_cell_out_Payload_in(36) [2]), .I (
         \uni_cell_out_Payload_in(36)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(36)(3)  (.O (
         \uni_cell_out_Payload_in(36) [3]), .I (
         \uni_cell_out_Payload_in(36)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(36)(4)  (.O (
         \uni_cell_out_Payload_in(36) [4]), .I (
         \uni_cell_out_Payload_in(36)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(36)(5)  (.O (
         \uni_cell_out_Payload_in(36) [5]), .I (
         \uni_cell_out_Payload_in(36)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(36)(6)  (.O (
         \uni_cell_out_Payload_in(36) [6]), .I (
         \uni_cell_out_Payload_in(36)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(36)(7)  (.O (
         \uni_cell_out_Payload_in(36) [7]), .I (
         \uni_cell_out_Payload_in(36)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(37)(0)  (.O (
         \uni_cell_out_Payload_in(37) [0]), .I (
         \uni_cell_out_Payload_in(37)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(37)(1)  (.O (
         \uni_cell_out_Payload_in(37) [1]), .I (
         \uni_cell_out_Payload_in(37)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(37)(2)  (.O (
         \uni_cell_out_Payload_in(37) [2]), .I (
         \uni_cell_out_Payload_in(37)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(37)(3)  (.O (
         \uni_cell_out_Payload_in(37) [3]), .I (
         \uni_cell_out_Payload_in(37)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(37)(4)  (.O (
         \uni_cell_out_Payload_in(37) [4]), .I (
         \uni_cell_out_Payload_in(37)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(37)(5)  (.O (
         \uni_cell_out_Payload_in(37) [5]), .I (
         \uni_cell_out_Payload_in(37)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(37)(6)  (.O (
         \uni_cell_out_Payload_in(37) [6]), .I (
         \uni_cell_out_Payload_in(37)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(37)(7)  (.O (
         \uni_cell_out_Payload_in(37) [7]), .I (
         \uni_cell_out_Payload_in(37)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(38)(0)  (.O (
         \uni_cell_out_Payload_in(38) [0]), .I (
         \uni_cell_out_Payload_in(38)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(38)(1)  (.O (
         \uni_cell_out_Payload_in(38) [1]), .I (
         \uni_cell_out_Payload_in(38)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(38)(2)  (.O (
         \uni_cell_out_Payload_in(38) [2]), .I (
         \uni_cell_out_Payload_in(38)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(38)(3)  (.O (
         \uni_cell_out_Payload_in(38) [3]), .I (
         \uni_cell_out_Payload_in(38)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(38)(4)  (.O (
         \uni_cell_out_Payload_in(38) [4]), .I (
         \uni_cell_out_Payload_in(38)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(38)(5)  (.O (
         \uni_cell_out_Payload_in(38) [5]), .I (
         \uni_cell_out_Payload_in(38)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(38)(6)  (.O (
         \uni_cell_out_Payload_in(38) [6]), .I (
         \uni_cell_out_Payload_in(38)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(38)(7)  (.O (
         \uni_cell_out_Payload_in(38) [7]), .I (
         \uni_cell_out_Payload_in(38)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(39)(0)  (.O (
         \uni_cell_out_Payload_in(39) [0]), .I (
         \uni_cell_out_Payload_in(39)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(39)(1)  (.O (
         \uni_cell_out_Payload_in(39) [1]), .I (
         \uni_cell_out_Payload_in(39)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(39)(2)  (.O (
         \uni_cell_out_Payload_in(39) [2]), .I (
         \uni_cell_out_Payload_in(39)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(39)(3)  (.O (
         \uni_cell_out_Payload_in(39) [3]), .I (
         \uni_cell_out_Payload_in(39)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(39)(4)  (.O (
         \uni_cell_out_Payload_in(39) [4]), .I (
         \uni_cell_out_Payload_in(39)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(39)(5)  (.O (
         \uni_cell_out_Payload_in(39) [5]), .I (
         \uni_cell_out_Payload_in(39)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(39)(6)  (.O (
         \uni_cell_out_Payload_in(39) [6]), .I (
         \uni_cell_out_Payload_in(39)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(39)(7)  (.O (
         \uni_cell_out_Payload_in(39) [7]), .I (
         \uni_cell_out_Payload_in(39)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(40)(0)  (.O (
         \uni_cell_out_Payload_in(40) [0]), .I (
         \uni_cell_out_Payload_in(40)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(40)(1)  (.O (
         \uni_cell_out_Payload_in(40) [1]), .I (
         \uni_cell_out_Payload_in(40)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(40)(2)  (.O (
         \uni_cell_out_Payload_in(40) [2]), .I (
         \uni_cell_out_Payload_in(40)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(40)(3)  (.O (
         \uni_cell_out_Payload_in(40) [3]), .I (
         \uni_cell_out_Payload_in(40)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(40)(4)  (.O (
         \uni_cell_out_Payload_in(40) [4]), .I (
         \uni_cell_out_Payload_in(40)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(40)(5)  (.O (
         \uni_cell_out_Payload_in(40) [5]), .I (
         \uni_cell_out_Payload_in(40)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(40)(6)  (.O (
         \uni_cell_out_Payload_in(40) [6]), .I (
         \uni_cell_out_Payload_in(40)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(40)(7)  (.O (
         \uni_cell_out_Payload_in(40) [7]), .I (
         \uni_cell_out_Payload_in(40)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(41)(0)  (.O (
         \uni_cell_out_Payload_in(41) [0]), .I (
         \uni_cell_out_Payload_in(41)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(41)(1)  (.O (
         \uni_cell_out_Payload_in(41) [1]), .I (
         \uni_cell_out_Payload_in(41)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(41)(2)  (.O (
         \uni_cell_out_Payload_in(41) [2]), .I (
         \uni_cell_out_Payload_in(41)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(41)(3)  (.O (
         \uni_cell_out_Payload_in(41) [3]), .I (
         \uni_cell_out_Payload_in(41)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(41)(4)  (.O (
         \uni_cell_out_Payload_in(41) [4]), .I (
         \uni_cell_out_Payload_in(41)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(41)(5)  (.O (
         \uni_cell_out_Payload_in(41) [5]), .I (
         \uni_cell_out_Payload_in(41)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(41)(6)  (.O (
         \uni_cell_out_Payload_in(41) [6]), .I (
         \uni_cell_out_Payload_in(41)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(41)(7)  (.O (
         \uni_cell_out_Payload_in(41) [7]), .I (
         \uni_cell_out_Payload_in(41)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(42)(0)  (.O (
         \uni_cell_out_Payload_in(42) [0]), .I (
         \uni_cell_out_Payload_in(42)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(42)(1)  (.O (
         \uni_cell_out_Payload_in(42) [1]), .I (
         \uni_cell_out_Payload_in(42)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(42)(2)  (.O (
         \uni_cell_out_Payload_in(42) [2]), .I (
         \uni_cell_out_Payload_in(42)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(42)(3)  (.O (
         \uni_cell_out_Payload_in(42) [3]), .I (
         \uni_cell_out_Payload_in(42)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(42)(4)  (.O (
         \uni_cell_out_Payload_in(42) [4]), .I (
         \uni_cell_out_Payload_in(42)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(42)(5)  (.O (
         \uni_cell_out_Payload_in(42) [5]), .I (
         \uni_cell_out_Payload_in(42)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(42)(6)  (.O (
         \uni_cell_out_Payload_in(42) [6]), .I (
         \uni_cell_out_Payload_in(42)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(42)(7)  (.O (
         \uni_cell_out_Payload_in(42) [7]), .I (
         \uni_cell_out_Payload_in(42)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(43)(0)  (.O (
         \uni_cell_out_Payload_in(43) [0]), .I (
         \uni_cell_out_Payload_in(43)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(43)(1)  (.O (
         \uni_cell_out_Payload_in(43) [1]), .I (
         \uni_cell_out_Payload_in(43)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(43)(2)  (.O (
         \uni_cell_out_Payload_in(43) [2]), .I (
         \uni_cell_out_Payload_in(43)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(43)(3)  (.O (
         \uni_cell_out_Payload_in(43) [3]), .I (
         \uni_cell_out_Payload_in(43)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(43)(4)  (.O (
         \uni_cell_out_Payload_in(43) [4]), .I (
         \uni_cell_out_Payload_in(43)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(43)(5)  (.O (
         \uni_cell_out_Payload_in(43) [5]), .I (
         \uni_cell_out_Payload_in(43)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(43)(6)  (.O (
         \uni_cell_out_Payload_in(43) [6]), .I (
         \uni_cell_out_Payload_in(43)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(43)(7)  (.O (
         \uni_cell_out_Payload_in(43) [7]), .I (
         \uni_cell_out_Payload_in(43)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(44)(0)  (.O (
         \uni_cell_out_Payload_in(44) [0]), .I (
         \uni_cell_out_Payload_in(44)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(44)(1)  (.O (
         \uni_cell_out_Payload_in(44) [1]), .I (
         \uni_cell_out_Payload_in(44)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(44)(2)  (.O (
         \uni_cell_out_Payload_in(44) [2]), .I (
         \uni_cell_out_Payload_in(44)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(44)(3)  (.O (
         \uni_cell_out_Payload_in(44) [3]), .I (
         \uni_cell_out_Payload_in(44)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(44)(4)  (.O (
         \uni_cell_out_Payload_in(44) [4]), .I (
         \uni_cell_out_Payload_in(44)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(44)(5)  (.O (
         \uni_cell_out_Payload_in(44) [5]), .I (
         \uni_cell_out_Payload_in(44)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(44)(6)  (.O (
         \uni_cell_out_Payload_in(44) [6]), .I (
         \uni_cell_out_Payload_in(44)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(44)(7)  (.O (
         \uni_cell_out_Payload_in(44) [7]), .I (
         \uni_cell_out_Payload_in(44)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(45)(0)  (.O (
         \uni_cell_out_Payload_in(45) [0]), .I (
         \uni_cell_out_Payload_in(45)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(45)(1)  (.O (
         \uni_cell_out_Payload_in(45) [1]), .I (
         \uni_cell_out_Payload_in(45)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(45)(2)  (.O (
         \uni_cell_out_Payload_in(45) [2]), .I (
         \uni_cell_out_Payload_in(45)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(45)(3)  (.O (
         \uni_cell_out_Payload_in(45) [3]), .I (
         \uni_cell_out_Payload_in(45)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(45)(4)  (.O (
         \uni_cell_out_Payload_in(45) [4]), .I (
         \uni_cell_out_Payload_in(45)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(45)(5)  (.O (
         \uni_cell_out_Payload_in(45) [5]), .I (
         \uni_cell_out_Payload_in(45)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(45)(6)  (.O (
         \uni_cell_out_Payload_in(45) [6]), .I (
         \uni_cell_out_Payload_in(45)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(45)(7)  (.O (
         \uni_cell_out_Payload_in(45) [7]), .I (
         \uni_cell_out_Payload_in(45)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(46)(0)  (.O (
         \uni_cell_out_Payload_in(46) [0]), .I (
         \uni_cell_out_Payload_in(46)_dup_0(0)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(46)(1)  (.O (
         \uni_cell_out_Payload_in(46) [1]), .I (
         \uni_cell_out_Payload_in(46)_dup_0(1)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(46)(2)  (.O (
         \uni_cell_out_Payload_in(46) [2]), .I (
         \uni_cell_out_Payload_in(46)_dup_0(2)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(46)(3)  (.O (
         \uni_cell_out_Payload_in(46) [3]), .I (
         \uni_cell_out_Payload_in(46)_dup_0(3)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(46)(4)  (.O (
         \uni_cell_out_Payload_in(46) [4]), .I (
         \uni_cell_out_Payload_in(46)_dup_0(4)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(46)(5)  (.O (
         \uni_cell_out_Payload_in(46) [5]), .I (
         \uni_cell_out_Payload_in(46)_dup_0(5)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(46)(6)  (.O (
         \uni_cell_out_Payload_in(46) [6]), .I (
         \uni_cell_out_Payload_in(46)_dup_0(6)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(46)(7)  (.O (
         \uni_cell_out_Payload_in(46) [7]), .I (
         \uni_cell_out_Payload_in(46)_dup_0(7)  )) ;
    OBUF \uni_cell_out_Payload_in_obuf(47)(0)  (.O (
         \uni_cell_out_Payload_in(47) [0]), .I (uni_cell_out_Payload_in_dup_0[0]
         )) ;
    OBUF \uni_cell_out_Payload_in_obuf(47)(1)  (.O (
         \uni_cell_out_Payload_in(47) [1]), .I (uni_cell_out_Payload_in_dup_0[1]
         )) ;
    OBUF \uni_cell_out_Payload_in_obuf(47)(2)  (.O (
         \uni_cell_out_Payload_in(47) [2]), .I (uni_cell_out_Payload_in_dup_0[2]
         )) ;
    OBUF \uni_cell_out_Payload_in_obuf(47)(3)  (.O (
         \uni_cell_out_Payload_in(47) [3]), .I (uni_cell_out_Payload_in_dup_0[3]
         )) ;
    OBUF \uni_cell_out_Payload_in_obuf(47)(4)  (.O (
         \uni_cell_out_Payload_in(47) [4]), .I (uni_cell_out_Payload_in_dup_0[4]
         )) ;
    OBUF \uni_cell_out_Payload_in_obuf(47)(5)  (.O (
         \uni_cell_out_Payload_in(47) [5]), .I (uni_cell_out_Payload_in_dup_0[5]
         )) ;
    OBUF \uni_cell_out_Payload_in_obuf(47)(6)  (.O (
         \uni_cell_out_Payload_in(47) [6]), .I (uni_cell_out_Payload_in_dup_0[6]
         )) ;
    OBUF \uni_cell_out_Payload_in_obuf(47)(7)  (.O (
         \uni_cell_out_Payload_in(47) [7]), .I (uni_cell_out_Payload_in_dup_0[7]
         )) ;
    IBUF \uni_cell_in_ibuf(0)  (.O (uni_cell_in_int[0]), .I (uni_cell_in[0])) ;
    IBUF \uni_cell_in_ibuf(1)  (.O (uni_cell_in_int[1]), .I (uni_cell_in[1])) ;
    IBUF \uni_cell_in_ibuf(2)  (.O (uni_cell_in_int[2]), .I (uni_cell_in[2])) ;
    IBUF \uni_cell_in_ibuf(3)  (.O (uni_cell_in_int[3]), .I (uni_cell_in[3])) ;
    IBUF \uni_cell_in_ibuf(4)  (.O (uni_cell_in_int[4]), .I (uni_cell_in[4])) ;
    IBUF \uni_cell_in_ibuf(5)  (.O (uni_cell_in_int[5]), .I (uni_cell_in[5])) ;
    IBUF \uni_cell_in_ibuf(6)  (.O (uni_cell_in_int[6]), .I (uni_cell_in[6])) ;
    IBUF \uni_cell_in_ibuf(7)  (.O (uni_cell_in_int[7]), .I (uni_cell_in[7])) ;
    IBUF \uni_cell_in_ibuf(8)  (.O (uni_cell_in_int[8]), .I (uni_cell_in[8])) ;
    IBUF \uni_cell_in_ibuf(9)  (.O (uni_cell_in_int[9]), .I (uni_cell_in[9])) ;
    IBUF \uni_cell_in_ibuf(10)  (.O (uni_cell_in_int[10]), .I (uni_cell_in[10])
         ) ;
    IBUF \uni_cell_in_ibuf(11)  (.O (uni_cell_in_int[11]), .I (uni_cell_in[11])
         ) ;
    IBUF \uni_cell_in_ibuf(12)  (.O (uni_cell_in_int[12]), .I (uni_cell_in[12])
         ) ;
    IBUF \uni_cell_in_ibuf(13)  (.O (uni_cell_in_int[13]), .I (uni_cell_in[13])
         ) ;
    IBUF \uni_cell_in_ibuf(14)  (.O (uni_cell_in_int[14]), .I (uni_cell_in[14])
         ) ;
    IBUF \uni_cell_in_ibuf(15)  (.O (uni_cell_in_int[15]), .I (uni_cell_in[15])
         ) ;
    IBUF \uni_cell_in_ibuf(16)  (.O (uni_cell_in_int[16]), .I (uni_cell_in[16])
         ) ;
    IBUF \uni_cell_in_ibuf(17)  (.O (uni_cell_in_int[17]), .I (uni_cell_in[17])
         ) ;
    IBUF \uni_cell_in_ibuf(18)  (.O (uni_cell_in_int[18]), .I (uni_cell_in[18])
         ) ;
    IBUF \uni_cell_in_ibuf(19)  (.O (uni_cell_in_int[19]), .I (uni_cell_in[19])
         ) ;
    IBUF \uni_cell_in_ibuf(20)  (.O (uni_cell_in_int[20]), .I (uni_cell_in[20])
         ) ;
    IBUF \uni_cell_in_ibuf(21)  (.O (uni_cell_in_int[21]), .I (uni_cell_in[21])
         ) ;
    IBUF \uni_cell_in_ibuf(22)  (.O (uni_cell_in_int[22]), .I (uni_cell_in[22])
         ) ;
    IBUF \uni_cell_in_ibuf(23)  (.O (uni_cell_in_int[23]), .I (uni_cell_in[23])
         ) ;
    IBUF \uni_cell_in_ibuf(24)  (.O (uni_cell_in_int[24]), .I (uni_cell_in[24])
         ) ;
    IBUF \uni_cell_in_ibuf(25)  (.O (uni_cell_in_int[25]), .I (uni_cell_in[25])
         ) ;
    IBUF \uni_cell_in_ibuf(26)  (.O (uni_cell_in_int[26]), .I (uni_cell_in[26])
         ) ;
    IBUF \uni_cell_in_ibuf(27)  (.O (uni_cell_in_int[27]), .I (uni_cell_in[27])
         ) ;
    IBUF \uni_cell_in_ibuf(28)  (.O (uni_cell_in_int[28]), .I (uni_cell_in[28])
         ) ;
    IBUF \uni_cell_in_ibuf(29)  (.O (uni_cell_in_int[29]), .I (uni_cell_in[29])
         ) ;
    IBUF \uni_cell_in_ibuf(30)  (.O (uni_cell_in_int[30]), .I (uni_cell_in[30])
         ) ;
    IBUF \uni_cell_in_ibuf(31)  (.O (uni_cell_in_int[31]), .I (uni_cell_in[31])
         ) ;
    IBUF \uni_cell_in_ibuf(32)  (.O (uni_cell_in_int[32]), .I (uni_cell_in[32])
         ) ;
    IBUF \uni_cell_in_ibuf(33)  (.O (uni_cell_in_int[33]), .I (uni_cell_in[33])
         ) ;
    IBUF \uni_cell_in_ibuf(34)  (.O (uni_cell_in_int[34]), .I (uni_cell_in[34])
         ) ;
    IBUF \uni_cell_in_ibuf(35)  (.O (uni_cell_in_int[35]), .I (uni_cell_in[35])
         ) ;
    IBUF \uni_cell_in_ibuf(36)  (.O (uni_cell_in_int[36]), .I (uni_cell_in[36])
         ) ;
    IBUF \uni_cell_in_ibuf(37)  (.O (uni_cell_in_int[37]), .I (uni_cell_in[37])
         ) ;
    IBUF \uni_cell_in_ibuf(38)  (.O (uni_cell_in_int[38]), .I (uni_cell_in[38])
         ) ;
    IBUF \uni_cell_in_ibuf(39)  (.O (uni_cell_in_int[39]), .I (uni_cell_in[39])
         ) ;
    IBUF \uni_cell_in_ibuf(40)  (.O (uni_cell_in_int[40]), .I (uni_cell_in[40])
         ) ;
    IBUF \uni_cell_in_ibuf(41)  (.O (uni_cell_in_int[41]), .I (uni_cell_in[41])
         ) ;
    IBUF \uni_cell_in_ibuf(42)  (.O (uni_cell_in_int[42]), .I (uni_cell_in[42])
         ) ;
    IBUF \uni_cell_in_ibuf(43)  (.O (uni_cell_in_int[43]), .I (uni_cell_in[43])
         ) ;
    IBUF \uni_cell_in_ibuf(44)  (.O (uni_cell_in_int[44]), .I (uni_cell_in[44])
         ) ;
    IBUF \uni_cell_in_ibuf(45)  (.O (uni_cell_in_int[45]), .I (uni_cell_in[45])
         ) ;
    IBUF \uni_cell_in_ibuf(46)  (.O (uni_cell_in_int[46]), .I (uni_cell_in[46])
         ) ;
    IBUF \uni_cell_in_ibuf(47)  (.O (uni_cell_in_int[47]), .I (uni_cell_in[47])
         ) ;
    IBUF \uni_cell_in_ibuf(48)  (.O (uni_cell_in_int[48]), .I (uni_cell_in[48])
         ) ;
    IBUF \uni_cell_in_ibuf(49)  (.O (uni_cell_in_int[49]), .I (uni_cell_in[49])
         ) ;
    IBUF \uni_cell_in_ibuf(50)  (.O (uni_cell_in_int[50]), .I (uni_cell_in[50])
         ) ;
    IBUF \uni_cell_in_ibuf(51)  (.O (uni_cell_in_int[51]), .I (uni_cell_in[51])
         ) ;
    IBUF \uni_cell_in_ibuf(52)  (.O (uni_cell_in_int[52]), .I (uni_cell_in[52])
         ) ;
    IBUF \uni_cell_in_ibuf(53)  (.O (uni_cell_in_int[53]), .I (uni_cell_in[53])
         ) ;
    IBUF \uni_cell_in_ibuf(54)  (.O (uni_cell_in_int[54]), .I (uni_cell_in[54])
         ) ;
    IBUF \uni_cell_in_ibuf(55)  (.O (uni_cell_in_int[55]), .I (uni_cell_in[55])
         ) ;
    IBUF \uni_cell_in_ibuf(56)  (.O (uni_cell_in_int[56]), .I (uni_cell_in[56])
         ) ;
    IBUF \uni_cell_in_ibuf(57)  (.O (uni_cell_in_int[57]), .I (uni_cell_in[57])
         ) ;
    IBUF \uni_cell_in_ibuf(58)  (.O (uni_cell_in_int[58]), .I (uni_cell_in[58])
         ) ;
    IBUF \uni_cell_in_ibuf(59)  (.O (uni_cell_in_int[59]), .I (uni_cell_in[59])
         ) ;
    IBUF \uni_cell_in_ibuf(60)  (.O (uni_cell_in_int[60]), .I (uni_cell_in[60])
         ) ;
    IBUF \uni_cell_in_ibuf(61)  (.O (uni_cell_in_int[61]), .I (uni_cell_in[61])
         ) ;
    IBUF \uni_cell_in_ibuf(62)  (.O (uni_cell_in_int[62]), .I (uni_cell_in[62])
         ) ;
    IBUF \uni_cell_in_ibuf(63)  (.O (uni_cell_in_int[63]), .I (uni_cell_in[63])
         ) ;
    IBUF \uni_cell_in_ibuf(64)  (.O (uni_cell_in_int[64]), .I (uni_cell_in[64])
         ) ;
    IBUF \uni_cell_in_ibuf(65)  (.O (uni_cell_in_int[65]), .I (uni_cell_in[65])
         ) ;
    IBUF \uni_cell_in_ibuf(66)  (.O (uni_cell_in_int[66]), .I (uni_cell_in[66])
         ) ;
    IBUF \uni_cell_in_ibuf(67)  (.O (uni_cell_in_int[67]), .I (uni_cell_in[67])
         ) ;
    IBUF \uni_cell_in_ibuf(68)  (.O (uni_cell_in_int[68]), .I (uni_cell_in[68])
         ) ;
    IBUF \uni_cell_in_ibuf(69)  (.O (uni_cell_in_int[69]), .I (uni_cell_in[69])
         ) ;
    IBUF \uni_cell_in_ibuf(70)  (.O (uni_cell_in_int[70]), .I (uni_cell_in[70])
         ) ;
    IBUF \uni_cell_in_ibuf(71)  (.O (uni_cell_in_int[71]), .I (uni_cell_in[71])
         ) ;
    IBUF \uni_cell_in_ibuf(72)  (.O (uni_cell_in_int[72]), .I (uni_cell_in[72])
         ) ;
    IBUF \uni_cell_in_ibuf(73)  (.O (uni_cell_in_int[73]), .I (uni_cell_in[73])
         ) ;
    IBUF \uni_cell_in_ibuf(74)  (.O (uni_cell_in_int[74]), .I (uni_cell_in[74])
         ) ;
    IBUF \uni_cell_in_ibuf(75)  (.O (uni_cell_in_int[75]), .I (uni_cell_in[75])
         ) ;
    IBUF \uni_cell_in_ibuf(76)  (.O (uni_cell_in_int[76]), .I (uni_cell_in[76])
         ) ;
    IBUF \uni_cell_in_ibuf(77)  (.O (uni_cell_in_int[77]), .I (uni_cell_in[77])
         ) ;
    IBUF \uni_cell_in_ibuf(78)  (.O (uni_cell_in_int[78]), .I (uni_cell_in[78])
         ) ;
    IBUF \uni_cell_in_ibuf(79)  (.O (uni_cell_in_int[79]), .I (uni_cell_in[79])
         ) ;
    IBUF \uni_cell_in_ibuf(80)  (.O (uni_cell_in_int[80]), .I (uni_cell_in[80])
         ) ;
    IBUF \uni_cell_in_ibuf(81)  (.O (uni_cell_in_int[81]), .I (uni_cell_in[81])
         ) ;
    IBUF \uni_cell_in_ibuf(82)  (.O (uni_cell_in_int[82]), .I (uni_cell_in[82])
         ) ;
    IBUF \uni_cell_in_ibuf(83)  (.O (uni_cell_in_int[83]), .I (uni_cell_in[83])
         ) ;
    IBUF \uni_cell_in_ibuf(84)  (.O (uni_cell_in_int[84]), .I (uni_cell_in[84])
         ) ;
    IBUF \uni_cell_in_ibuf(85)  (.O (uni_cell_in_int[85]), .I (uni_cell_in[85])
         ) ;
    IBUF \uni_cell_in_ibuf(86)  (.O (uni_cell_in_int[86]), .I (uni_cell_in[86])
         ) ;
    IBUF \uni_cell_in_ibuf(87)  (.O (uni_cell_in_int[87]), .I (uni_cell_in[87])
         ) ;
    IBUF \uni_cell_in_ibuf(88)  (.O (uni_cell_in_int[88]), .I (uni_cell_in[88])
         ) ;
    IBUF \uni_cell_in_ibuf(89)  (.O (uni_cell_in_int[89]), .I (uni_cell_in[89])
         ) ;
    IBUF \uni_cell_in_ibuf(90)  (.O (uni_cell_in_int[90]), .I (uni_cell_in[90])
         ) ;
    IBUF \uni_cell_in_ibuf(91)  (.O (uni_cell_in_int[91]), .I (uni_cell_in[91])
         ) ;
    IBUF \uni_cell_in_ibuf(92)  (.O (uni_cell_in_int[92]), .I (uni_cell_in[92])
         ) ;
    IBUF \uni_cell_in_ibuf(93)  (.O (uni_cell_in_int[93]), .I (uni_cell_in[93])
         ) ;
    IBUF \uni_cell_in_ibuf(94)  (.O (uni_cell_in_int[94]), .I (uni_cell_in[94])
         ) ;
    IBUF \uni_cell_in_ibuf(95)  (.O (uni_cell_in_int[95]), .I (uni_cell_in[95])
         ) ;
    IBUF \uni_cell_in_ibuf(96)  (.O (uni_cell_in_int[96]), .I (uni_cell_in[96])
         ) ;
    IBUF \uni_cell_in_ibuf(97)  (.O (uni_cell_in_int[97]), .I (uni_cell_in[97])
         ) ;
    IBUF \uni_cell_in_ibuf(98)  (.O (uni_cell_in_int[98]), .I (uni_cell_in[98])
         ) ;
    IBUF \uni_cell_in_ibuf(99)  (.O (uni_cell_in_int[99]), .I (uni_cell_in[99])
         ) ;
    IBUF \uni_cell_in_ibuf(100)  (.O (uni_cell_in_int[100]), .I (
         uni_cell_in[100])) ;
    IBUF \uni_cell_in_ibuf(101)  (.O (uni_cell_in_int[101]), .I (
         uni_cell_in[101])) ;
    IBUF \uni_cell_in_ibuf(102)  (.O (uni_cell_in_int[102]), .I (
         uni_cell_in[102])) ;
    IBUF \uni_cell_in_ibuf(103)  (.O (uni_cell_in_int[103]), .I (
         uni_cell_in[103])) ;
    IBUF \uni_cell_in_ibuf(104)  (.O (uni_cell_in_int[104]), .I (
         uni_cell_in[104])) ;
    IBUF \uni_cell_in_ibuf(105)  (.O (uni_cell_in_int[105]), .I (
         uni_cell_in[105])) ;
    IBUF \uni_cell_in_ibuf(106)  (.O (uni_cell_in_int[106]), .I (
         uni_cell_in[106])) ;
    IBUF \uni_cell_in_ibuf(107)  (.O (uni_cell_in_int[107]), .I (
         uni_cell_in[107])) ;
    IBUF \uni_cell_in_ibuf(108)  (.O (uni_cell_in_int[108]), .I (
         uni_cell_in[108])) ;
    IBUF \uni_cell_in_ibuf(109)  (.O (uni_cell_in_int[109]), .I (
         uni_cell_in[109])) ;
    IBUF \uni_cell_in_ibuf(110)  (.O (uni_cell_in_int[110]), .I (
         uni_cell_in[110])) ;
    IBUF \uni_cell_in_ibuf(111)  (.O (uni_cell_in_int[111]), .I (
         uni_cell_in[111])) ;
    IBUF \uni_cell_in_ibuf(112)  (.O (uni_cell_in_int[112]), .I (
         uni_cell_in[112])) ;
    IBUF \uni_cell_in_ibuf(113)  (.O (uni_cell_in_int[113]), .I (
         uni_cell_in[113])) ;
    IBUF \uni_cell_in_ibuf(114)  (.O (uni_cell_in_int[114]), .I (
         uni_cell_in[114])) ;
    IBUF \uni_cell_in_ibuf(115)  (.O (uni_cell_in_int[115]), .I (
         uni_cell_in[115])) ;
    IBUF \uni_cell_in_ibuf(116)  (.O (uni_cell_in_int[116]), .I (
         uni_cell_in[116])) ;
    IBUF \uni_cell_in_ibuf(117)  (.O (uni_cell_in_int[117]), .I (
         uni_cell_in[117])) ;
    IBUF \uni_cell_in_ibuf(118)  (.O (uni_cell_in_int[118]), .I (
         uni_cell_in[118])) ;
    IBUF \uni_cell_in_ibuf(119)  (.O (uni_cell_in_int[119]), .I (
         uni_cell_in[119])) ;
    IBUF \uni_cell_in_ibuf(120)  (.O (uni_cell_in_int[120]), .I (
         uni_cell_in[120])) ;
    IBUF \uni_cell_in_ibuf(121)  (.O (uni_cell_in_int[121]), .I (
         uni_cell_in[121])) ;
    IBUF \uni_cell_in_ibuf(122)  (.O (uni_cell_in_int[122]), .I (
         uni_cell_in[122])) ;
    IBUF \uni_cell_in_ibuf(123)  (.O (uni_cell_in_int[123]), .I (
         uni_cell_in[123])) ;
    IBUF \uni_cell_in_ibuf(124)  (.O (uni_cell_in_int[124]), .I (
         uni_cell_in[124])) ;
    IBUF \uni_cell_in_ibuf(125)  (.O (uni_cell_in_int[125]), .I (
         uni_cell_in[125])) ;
    IBUF \uni_cell_in_ibuf(126)  (.O (uni_cell_in_int[126]), .I (
         uni_cell_in[126])) ;
    IBUF \uni_cell_in_ibuf(127)  (.O (uni_cell_in_int[127]), .I (
         uni_cell_in[127])) ;
    IBUF \uni_cell_in_ibuf(128)  (.O (uni_cell_in_int[128]), .I (
         uni_cell_in[128])) ;
    IBUF \uni_cell_in_ibuf(129)  (.O (uni_cell_in_int[129]), .I (
         uni_cell_in[129])) ;
    IBUF \uni_cell_in_ibuf(130)  (.O (uni_cell_in_int[130]), .I (
         uni_cell_in[130])) ;
    IBUF \uni_cell_in_ibuf(131)  (.O (uni_cell_in_int[131]), .I (
         uni_cell_in[131])) ;
    IBUF \uni_cell_in_ibuf(132)  (.O (uni_cell_in_int[132]), .I (
         uni_cell_in[132])) ;
    IBUF \uni_cell_in_ibuf(133)  (.O (uni_cell_in_int[133]), .I (
         uni_cell_in[133])) ;
    IBUF \uni_cell_in_ibuf(134)  (.O (uni_cell_in_int[134]), .I (
         uni_cell_in[134])) ;
    IBUF \uni_cell_in_ibuf(135)  (.O (uni_cell_in_int[135]), .I (
         uni_cell_in[135])) ;
    IBUF \uni_cell_in_ibuf(136)  (.O (uni_cell_in_int[136]), .I (
         uni_cell_in[136])) ;
    IBUF \uni_cell_in_ibuf(137)  (.O (uni_cell_in_int[137]), .I (
         uni_cell_in[137])) ;
    IBUF \uni_cell_in_ibuf(138)  (.O (uni_cell_in_int[138]), .I (
         uni_cell_in[138])) ;
    IBUF \uni_cell_in_ibuf(139)  (.O (uni_cell_in_int[139]), .I (
         uni_cell_in[139])) ;
    IBUF \uni_cell_in_ibuf(140)  (.O (uni_cell_in_int[140]), .I (
         uni_cell_in[140])) ;
    IBUF \uni_cell_in_ibuf(141)  (.O (uni_cell_in_int[141]), .I (
         uni_cell_in[141])) ;
    IBUF \uni_cell_in_ibuf(142)  (.O (uni_cell_in_int[142]), .I (
         uni_cell_in[142])) ;
    IBUF \uni_cell_in_ibuf(143)  (.O (uni_cell_in_int[143]), .I (
         uni_cell_in[143])) ;
    IBUF \uni_cell_in_ibuf(144)  (.O (uni_cell_in_int[144]), .I (
         uni_cell_in[144])) ;
    IBUF \uni_cell_in_ibuf(145)  (.O (uni_cell_in_int[145]), .I (
         uni_cell_in[145])) ;
    IBUF \uni_cell_in_ibuf(146)  (.O (uni_cell_in_int[146]), .I (
         uni_cell_in[146])) ;
    IBUF \uni_cell_in_ibuf(147)  (.O (uni_cell_in_int[147]), .I (
         uni_cell_in[147])) ;
    IBUF \uni_cell_in_ibuf(148)  (.O (uni_cell_in_int[148]), .I (
         uni_cell_in[148])) ;
    IBUF \uni_cell_in_ibuf(149)  (.O (uni_cell_in_int[149]), .I (
         uni_cell_in[149])) ;
    IBUF \uni_cell_in_ibuf(150)  (.O (uni_cell_in_int[150]), .I (
         uni_cell_in[150])) ;
    IBUF \uni_cell_in_ibuf(151)  (.O (uni_cell_in_int[151]), .I (
         uni_cell_in[151])) ;
    IBUF \uni_cell_in_ibuf(152)  (.O (uni_cell_in_int[152]), .I (
         uni_cell_in[152])) ;
    IBUF \uni_cell_in_ibuf(153)  (.O (uni_cell_in_int[153]), .I (
         uni_cell_in[153])) ;
    IBUF \uni_cell_in_ibuf(154)  (.O (uni_cell_in_int[154]), .I (
         uni_cell_in[154])) ;
    IBUF \uni_cell_in_ibuf(155)  (.O (uni_cell_in_int[155]), .I (
         uni_cell_in[155])) ;
    IBUF \uni_cell_in_ibuf(156)  (.O (uni_cell_in_int[156]), .I (
         uni_cell_in[156])) ;
    IBUF \uni_cell_in_ibuf(157)  (.O (uni_cell_in_int[157]), .I (
         uni_cell_in[157])) ;
    IBUF \uni_cell_in_ibuf(158)  (.O (uni_cell_in_int[158]), .I (
         uni_cell_in[158])) ;
    IBUF \uni_cell_in_ibuf(159)  (.O (uni_cell_in_int[159]), .I (
         uni_cell_in[159])) ;
    IBUF \uni_cell_in_ibuf(160)  (.O (uni_cell_in_int[160]), .I (
         uni_cell_in[160])) ;
    IBUF \uni_cell_in_ibuf(161)  (.O (uni_cell_in_int[161]), .I (
         uni_cell_in[161])) ;
    IBUF \uni_cell_in_ibuf(162)  (.O (uni_cell_in_int[162]), .I (
         uni_cell_in[162])) ;
    IBUF \uni_cell_in_ibuf(163)  (.O (uni_cell_in_int[163]), .I (
         uni_cell_in[163])) ;
    IBUF \uni_cell_in_ibuf(164)  (.O (uni_cell_in_int[164]), .I (
         uni_cell_in[164])) ;
    IBUF \uni_cell_in_ibuf(165)  (.O (uni_cell_in_int[165]), .I (
         uni_cell_in[165])) ;
    IBUF \uni_cell_in_ibuf(166)  (.O (uni_cell_in_int[166]), .I (
         uni_cell_in[166])) ;
    IBUF \uni_cell_in_ibuf(167)  (.O (uni_cell_in_int[167]), .I (
         uni_cell_in[167])) ;
    IBUF \uni_cell_in_ibuf(168)  (.O (uni_cell_in_int[168]), .I (
         uni_cell_in[168])) ;
    IBUF \uni_cell_in_ibuf(169)  (.O (uni_cell_in_int[169]), .I (
         uni_cell_in[169])) ;
    IBUF \uni_cell_in_ibuf(170)  (.O (uni_cell_in_int[170]), .I (
         uni_cell_in[170])) ;
    IBUF \uni_cell_in_ibuf(171)  (.O (uni_cell_in_int[171]), .I (
         uni_cell_in[171])) ;
    IBUF \uni_cell_in_ibuf(172)  (.O (uni_cell_in_int[172]), .I (
         uni_cell_in[172])) ;
    IBUF \uni_cell_in_ibuf(173)  (.O (uni_cell_in_int[173]), .I (
         uni_cell_in[173])) ;
    IBUF \uni_cell_in_ibuf(174)  (.O (uni_cell_in_int[174]), .I (
         uni_cell_in[174])) ;
    IBUF \uni_cell_in_ibuf(175)  (.O (uni_cell_in_int[175]), .I (
         uni_cell_in[175])) ;
    IBUF \uni_cell_in_ibuf(176)  (.O (uni_cell_in_int[176]), .I (
         uni_cell_in[176])) ;
    IBUF \uni_cell_in_ibuf(177)  (.O (uni_cell_in_int[177]), .I (
         uni_cell_in[177])) ;
    IBUF \uni_cell_in_ibuf(178)  (.O (uni_cell_in_int[178]), .I (
         uni_cell_in[178])) ;
    IBUF \uni_cell_in_ibuf(179)  (.O (uni_cell_in_int[179]), .I (
         uni_cell_in[179])) ;
    IBUF \uni_cell_in_ibuf(180)  (.O (uni_cell_in_int[180]), .I (
         uni_cell_in[180])) ;
    IBUF \uni_cell_in_ibuf(181)  (.O (uni_cell_in_int[181]), .I (
         uni_cell_in[181])) ;
    IBUF \uni_cell_in_ibuf(182)  (.O (uni_cell_in_int[182]), .I (
         uni_cell_in[182])) ;
    IBUF \uni_cell_in_ibuf(183)  (.O (uni_cell_in_int[183]), .I (
         uni_cell_in[183])) ;
    IBUF \uni_cell_in_ibuf(184)  (.O (uni_cell_in_int[184]), .I (
         uni_cell_in[184])) ;
    IBUF \uni_cell_in_ibuf(185)  (.O (uni_cell_in_int[185]), .I (
         uni_cell_in[185])) ;
    IBUF \uni_cell_in_ibuf(186)  (.O (uni_cell_in_int[186]), .I (
         uni_cell_in[186])) ;
    IBUF \uni_cell_in_ibuf(187)  (.O (uni_cell_in_int[187]), .I (
         uni_cell_in[187])) ;
    IBUF \uni_cell_in_ibuf(188)  (.O (uni_cell_in_int[188]), .I (
         uni_cell_in[188])) ;
    IBUF \uni_cell_in_ibuf(189)  (.O (uni_cell_in_int[189]), .I (
         uni_cell_in[189])) ;
    IBUF \uni_cell_in_ibuf(190)  (.O (uni_cell_in_int[190]), .I (
         uni_cell_in[190])) ;
    IBUF \uni_cell_in_ibuf(191)  (.O (uni_cell_in_int[191]), .I (
         uni_cell_in[191])) ;
    IBUF \uni_cell_in_ibuf(192)  (.O (uni_cell_in_int[192]), .I (
         uni_cell_in[192])) ;
    IBUF \uni_cell_in_ibuf(193)  (.O (uni_cell_in_int[193]), .I (
         uni_cell_in[193])) ;
    IBUF \uni_cell_in_ibuf(194)  (.O (uni_cell_in_int[194]), .I (
         uni_cell_in[194])) ;
    IBUF \uni_cell_in_ibuf(195)  (.O (uni_cell_in_int[195]), .I (
         uni_cell_in[195])) ;
    IBUF \uni_cell_in_ibuf(196)  (.O (uni_cell_in_int[196]), .I (
         uni_cell_in[196])) ;
    IBUF \uni_cell_in_ibuf(197)  (.O (uni_cell_in_int[197]), .I (
         uni_cell_in[197])) ;
    IBUF \uni_cell_in_ibuf(198)  (.O (uni_cell_in_int[198]), .I (
         uni_cell_in[198])) ;
    IBUF \uni_cell_in_ibuf(199)  (.O (uni_cell_in_int[199]), .I (
         uni_cell_in[199])) ;
    IBUF \uni_cell_in_ibuf(200)  (.O (uni_cell_in_int[200]), .I (
         uni_cell_in[200])) ;
    IBUF \uni_cell_in_ibuf(201)  (.O (uni_cell_in_int[201]), .I (
         uni_cell_in[201])) ;
    IBUF \uni_cell_in_ibuf(202)  (.O (uni_cell_in_int[202]), .I (
         uni_cell_in[202])) ;
    IBUF \uni_cell_in_ibuf(203)  (.O (uni_cell_in_int[203]), .I (
         uni_cell_in[203])) ;
    IBUF \uni_cell_in_ibuf(204)  (.O (uni_cell_in_int[204]), .I (
         uni_cell_in[204])) ;
    IBUF \uni_cell_in_ibuf(205)  (.O (uni_cell_in_int[205]), .I (
         uni_cell_in[205])) ;
    IBUF \uni_cell_in_ibuf(206)  (.O (uni_cell_in_int[206]), .I (
         uni_cell_in[206])) ;
    IBUF \uni_cell_in_ibuf(207)  (.O (uni_cell_in_int[207]), .I (
         uni_cell_in[207])) ;
    IBUF \uni_cell_in_ibuf(208)  (.O (uni_cell_in_int[208]), .I (
         uni_cell_in[208])) ;
    IBUF \uni_cell_in_ibuf(209)  (.O (uni_cell_in_int[209]), .I (
         uni_cell_in[209])) ;
    IBUF \uni_cell_in_ibuf(210)  (.O (uni_cell_in_int[210]), .I (
         uni_cell_in[210])) ;
    IBUF \uni_cell_in_ibuf(211)  (.O (uni_cell_in_int[211]), .I (
         uni_cell_in[211])) ;
    IBUF \uni_cell_in_ibuf(212)  (.O (uni_cell_in_int[212]), .I (
         uni_cell_in[212])) ;
    IBUF \uni_cell_in_ibuf(213)  (.O (uni_cell_in_int[213]), .I (
         uni_cell_in[213])) ;
    IBUF \uni_cell_in_ibuf(214)  (.O (uni_cell_in_int[214]), .I (
         uni_cell_in[214])) ;
    IBUF \uni_cell_in_ibuf(215)  (.O (uni_cell_in_int[215]), .I (
         uni_cell_in[215])) ;
    IBUF \uni_cell_in_ibuf(216)  (.O (uni_cell_in_int[216]), .I (
         uni_cell_in[216])) ;
    IBUF \uni_cell_in_ibuf(217)  (.O (uni_cell_in_int[217]), .I (
         uni_cell_in[217])) ;
    IBUF \uni_cell_in_ibuf(218)  (.O (uni_cell_in_int[218]), .I (
         uni_cell_in[218])) ;
    IBUF \uni_cell_in_ibuf(219)  (.O (uni_cell_in_int[219]), .I (
         uni_cell_in[219])) ;
    IBUF \uni_cell_in_ibuf(220)  (.O (uni_cell_in_int[220]), .I (
         uni_cell_in[220])) ;
    IBUF \uni_cell_in_ibuf(221)  (.O (uni_cell_in_int[221]), .I (
         uni_cell_in[221])) ;
    IBUF \uni_cell_in_ibuf(222)  (.O (uni_cell_in_int[222]), .I (
         uni_cell_in[222])) ;
    IBUF \uni_cell_in_ibuf(223)  (.O (uni_cell_in_int[223]), .I (
         uni_cell_in[223])) ;
    IBUF \uni_cell_in_ibuf(224)  (.O (uni_cell_in_int[224]), .I (
         uni_cell_in[224])) ;
    IBUF \uni_cell_in_ibuf(225)  (.O (uni_cell_in_int[225]), .I (
         uni_cell_in[225])) ;
    IBUF \uni_cell_in_ibuf(226)  (.O (uni_cell_in_int[226]), .I (
         uni_cell_in[226])) ;
    IBUF \uni_cell_in_ibuf(227)  (.O (uni_cell_in_int[227]), .I (
         uni_cell_in[227])) ;
    IBUF \uni_cell_in_ibuf(228)  (.O (uni_cell_in_int[228]), .I (
         uni_cell_in[228])) ;
    IBUF \uni_cell_in_ibuf(229)  (.O (uni_cell_in_int[229]), .I (
         uni_cell_in[229])) ;
    IBUF \uni_cell_in_ibuf(230)  (.O (uni_cell_in_int[230]), .I (
         uni_cell_in[230])) ;
    IBUF \uni_cell_in_ibuf(231)  (.O (uni_cell_in_int[231]), .I (
         uni_cell_in[231])) ;
    IBUF \uni_cell_in_ibuf(232)  (.O (uni_cell_in_int[232]), .I (
         uni_cell_in[232])) ;
    IBUF \uni_cell_in_ibuf(233)  (.O (uni_cell_in_int[233]), .I (
         uni_cell_in[233])) ;
    IBUF \uni_cell_in_ibuf(234)  (.O (uni_cell_in_int[234]), .I (
         uni_cell_in[234])) ;
    IBUF \uni_cell_in_ibuf(235)  (.O (uni_cell_in_int[235]), .I (
         uni_cell_in[235])) ;
    IBUF \uni_cell_in_ibuf(236)  (.O (uni_cell_in_int[236]), .I (
         uni_cell_in[236])) ;
    IBUF \uni_cell_in_ibuf(237)  (.O (uni_cell_in_int[237]), .I (
         uni_cell_in[237])) ;
    IBUF \uni_cell_in_ibuf(238)  (.O (uni_cell_in_int[238]), .I (
         uni_cell_in[238])) ;
    IBUF \uni_cell_in_ibuf(239)  (.O (uni_cell_in_int[239]), .I (
         uni_cell_in[239])) ;
    IBUF \uni_cell_in_ibuf(240)  (.O (uni_cell_in_int[240]), .I (
         uni_cell_in[240])) ;
    IBUF \uni_cell_in_ibuf(241)  (.O (uni_cell_in_int[241]), .I (
         uni_cell_in[241])) ;
    IBUF \uni_cell_in_ibuf(242)  (.O (uni_cell_in_int[242]), .I (
         uni_cell_in[242])) ;
    IBUF \uni_cell_in_ibuf(243)  (.O (uni_cell_in_int[243]), .I (
         uni_cell_in[243])) ;
    IBUF \uni_cell_in_ibuf(244)  (.O (uni_cell_in_int[244]), .I (
         uni_cell_in[244])) ;
    IBUF \uni_cell_in_ibuf(245)  (.O (uni_cell_in_int[245]), .I (
         uni_cell_in[245])) ;
    IBUF \uni_cell_in_ibuf(246)  (.O (uni_cell_in_int[246]), .I (
         uni_cell_in[246])) ;
    IBUF \uni_cell_in_ibuf(247)  (.O (uni_cell_in_int[247]), .I (
         uni_cell_in[247])) ;
    IBUF \uni_cell_in_ibuf(248)  (.O (uni_cell_in_int[248]), .I (
         uni_cell_in[248])) ;
    IBUF \uni_cell_in_ibuf(249)  (.O (uni_cell_in_int[249]), .I (
         uni_cell_in[249])) ;
    IBUF \uni_cell_in_ibuf(250)  (.O (uni_cell_in_int[250]), .I (
         uni_cell_in[250])) ;
    IBUF \uni_cell_in_ibuf(251)  (.O (uni_cell_in_int[251]), .I (
         uni_cell_in[251])) ;
    IBUF \uni_cell_in_ibuf(252)  (.O (uni_cell_in_int[252]), .I (
         uni_cell_in[252])) ;
    IBUF \uni_cell_in_ibuf(253)  (.O (uni_cell_in_int[253]), .I (
         uni_cell_in[253])) ;
    IBUF \uni_cell_in_ibuf(254)  (.O (uni_cell_in_int[254]), .I (
         uni_cell_in[254])) ;
    IBUF \uni_cell_in_ibuf(255)  (.O (uni_cell_in_int[255]), .I (
         uni_cell_in[255])) ;
    IBUF \uni_cell_in_ibuf(256)  (.O (uni_cell_in_int[256]), .I (
         uni_cell_in[256])) ;
    IBUF \uni_cell_in_ibuf(257)  (.O (uni_cell_in_int[257]), .I (
         uni_cell_in[257])) ;
    IBUF \uni_cell_in_ibuf(258)  (.O (uni_cell_in_int[258]), .I (
         uni_cell_in[258])) ;
    IBUF \uni_cell_in_ibuf(259)  (.O (uni_cell_in_int[259]), .I (
         uni_cell_in[259])) ;
    IBUF \uni_cell_in_ibuf(260)  (.O (uni_cell_in_int[260]), .I (
         uni_cell_in[260])) ;
    IBUF \uni_cell_in_ibuf(261)  (.O (uni_cell_in_int[261]), .I (
         uni_cell_in[261])) ;
    IBUF \uni_cell_in_ibuf(262)  (.O (uni_cell_in_int[262]), .I (
         uni_cell_in[262])) ;
    IBUF \uni_cell_in_ibuf(263)  (.O (uni_cell_in_int[263]), .I (
         uni_cell_in[263])) ;
    IBUF \uni_cell_in_ibuf(264)  (.O (uni_cell_in_int[264]), .I (
         uni_cell_in[264])) ;
    IBUF \uni_cell_in_ibuf(265)  (.O (uni_cell_in_int[265]), .I (
         uni_cell_in[265])) ;
    IBUF \uni_cell_in_ibuf(266)  (.O (uni_cell_in_int[266]), .I (
         uni_cell_in[266])) ;
    IBUF \uni_cell_in_ibuf(267)  (.O (uni_cell_in_int[267]), .I (
         uni_cell_in[267])) ;
    IBUF \uni_cell_in_ibuf(268)  (.O (uni_cell_in_int[268]), .I (
         uni_cell_in[268])) ;
    IBUF \uni_cell_in_ibuf(269)  (.O (uni_cell_in_int[269]), .I (
         uni_cell_in[269])) ;
    IBUF \uni_cell_in_ibuf(270)  (.O (uni_cell_in_int[270]), .I (
         uni_cell_in[270])) ;
    IBUF \uni_cell_in_ibuf(271)  (.O (uni_cell_in_int[271]), .I (
         uni_cell_in[271])) ;
    IBUF \uni_cell_in_ibuf(272)  (.O (uni_cell_in_int[272]), .I (
         uni_cell_in[272])) ;
    IBUF \uni_cell_in_ibuf(273)  (.O (uni_cell_in_int[273]), .I (
         uni_cell_in[273])) ;
    IBUF \uni_cell_in_ibuf(274)  (.O (uni_cell_in_int[274]), .I (
         uni_cell_in[274])) ;
    IBUF \uni_cell_in_ibuf(275)  (.O (uni_cell_in_int[275]), .I (
         uni_cell_in[275])) ;
    IBUF \uni_cell_in_ibuf(276)  (.O (uni_cell_in_int[276]), .I (
         uni_cell_in[276])) ;
    IBUF \uni_cell_in_ibuf(277)  (.O (uni_cell_in_int[277]), .I (
         uni_cell_in[277])) ;
    IBUF \uni_cell_in_ibuf(278)  (.O (uni_cell_in_int[278]), .I (
         uni_cell_in[278])) ;
    IBUF \uni_cell_in_ibuf(279)  (.O (uni_cell_in_int[279]), .I (
         uni_cell_in[279])) ;
    IBUF \uni_cell_in_ibuf(280)  (.O (uni_cell_in_int[280]), .I (
         uni_cell_in[280])) ;
    IBUF \uni_cell_in_ibuf(281)  (.O (uni_cell_in_int[281]), .I (
         uni_cell_in[281])) ;
    IBUF \uni_cell_in_ibuf(282)  (.O (uni_cell_in_int[282]), .I (
         uni_cell_in[282])) ;
    IBUF \uni_cell_in_ibuf(283)  (.O (uni_cell_in_int[283]), .I (
         uni_cell_in[283])) ;
    IBUF \uni_cell_in_ibuf(284)  (.O (uni_cell_in_int[284]), .I (
         uni_cell_in[284])) ;
    IBUF \uni_cell_in_ibuf(285)  (.O (uni_cell_in_int[285]), .I (
         uni_cell_in[285])) ;
    IBUF \uni_cell_in_ibuf(286)  (.O (uni_cell_in_int[286]), .I (
         uni_cell_in[286])) ;
    IBUF \uni_cell_in_ibuf(287)  (.O (uni_cell_in_int[287]), .I (
         uni_cell_in[287])) ;
    IBUF \uni_cell_in_ibuf(288)  (.O (uni_cell_in_int[288]), .I (
         uni_cell_in[288])) ;
    IBUF \uni_cell_in_ibuf(289)  (.O (uni_cell_in_int[289]), .I (
         uni_cell_in[289])) ;
    IBUF \uni_cell_in_ibuf(290)  (.O (uni_cell_in_int[290]), .I (
         uni_cell_in[290])) ;
    IBUF \uni_cell_in_ibuf(291)  (.O (uni_cell_in_int[291]), .I (
         uni_cell_in[291])) ;
    IBUF \uni_cell_in_ibuf(292)  (.O (uni_cell_in_int[292]), .I (
         uni_cell_in[292])) ;
    IBUF \uni_cell_in_ibuf(293)  (.O (uni_cell_in_int[293]), .I (
         uni_cell_in[293])) ;
    IBUF \uni_cell_in_ibuf(294)  (.O (uni_cell_in_int[294]), .I (
         uni_cell_in[294])) ;
    IBUF \uni_cell_in_ibuf(295)  (.O (uni_cell_in_int[295]), .I (
         uni_cell_in[295])) ;
    IBUF \uni_cell_in_ibuf(296)  (.O (uni_cell_in_int[296]), .I (
         uni_cell_in[296])) ;
    IBUF \uni_cell_in_ibuf(297)  (.O (uni_cell_in_int[297]), .I (
         uni_cell_in[297])) ;
    IBUF \uni_cell_in_ibuf(298)  (.O (uni_cell_in_int[298]), .I (
         uni_cell_in[298])) ;
    IBUF \uni_cell_in_ibuf(299)  (.O (uni_cell_in_int[299]), .I (
         uni_cell_in[299])) ;
    IBUF \uni_cell_in_ibuf(300)  (.O (uni_cell_in_int[300]), .I (
         uni_cell_in[300])) ;
    IBUF \uni_cell_in_ibuf(301)  (.O (uni_cell_in_int[301]), .I (
         uni_cell_in[301])) ;
    IBUF \uni_cell_in_ibuf(302)  (.O (uni_cell_in_int[302]), .I (
         uni_cell_in[302])) ;
    IBUF \uni_cell_in_ibuf(303)  (.O (uni_cell_in_int[303]), .I (
         uni_cell_in[303])) ;
    IBUF \uni_cell_in_ibuf(304)  (.O (uni_cell_in_int[304]), .I (
         uni_cell_in[304])) ;
    IBUF \uni_cell_in_ibuf(305)  (.O (uni_cell_in_int[305]), .I (
         uni_cell_in[305])) ;
    IBUF \uni_cell_in_ibuf(306)  (.O (uni_cell_in_int[306]), .I (
         uni_cell_in[306])) ;
    IBUF \uni_cell_in_ibuf(307)  (.O (uni_cell_in_int[307]), .I (
         uni_cell_in[307])) ;
    IBUF \uni_cell_in_ibuf(308)  (.O (uni_cell_in_int[308]), .I (
         uni_cell_in[308])) ;
    IBUF \uni_cell_in_ibuf(309)  (.O (uni_cell_in_int[309]), .I (
         uni_cell_in[309])) ;
    IBUF \uni_cell_in_ibuf(310)  (.O (uni_cell_in_int[310]), .I (
         uni_cell_in[310])) ;
    IBUF \uni_cell_in_ibuf(311)  (.O (uni_cell_in_int[311]), .I (
         uni_cell_in[311])) ;
    IBUF \uni_cell_in_ibuf(312)  (.O (uni_cell_in_int[312]), .I (
         uni_cell_in[312])) ;
    IBUF \uni_cell_in_ibuf(313)  (.O (uni_cell_in_int[313]), .I (
         uni_cell_in[313])) ;
    IBUF \uni_cell_in_ibuf(314)  (.O (uni_cell_in_int[314]), .I (
         uni_cell_in[314])) ;
    IBUF \uni_cell_in_ibuf(315)  (.O (uni_cell_in_int[315]), .I (
         uni_cell_in[315])) ;
    IBUF \uni_cell_in_ibuf(316)  (.O (uni_cell_in_int[316]), .I (
         uni_cell_in[316])) ;
    IBUF \uni_cell_in_ibuf(317)  (.O (uni_cell_in_int[317]), .I (
         uni_cell_in[317])) ;
    IBUF \uni_cell_in_ibuf(318)  (.O (uni_cell_in_int[318]), .I (
         uni_cell_in[318])) ;
    IBUF \uni_cell_in_ibuf(319)  (.O (uni_cell_in_int[319]), .I (
         uni_cell_in[319])) ;
    IBUF \uni_cell_in_ibuf(320)  (.O (uni_cell_in_int[320]), .I (
         uni_cell_in[320])) ;
    IBUF \uni_cell_in_ibuf(321)  (.O (uni_cell_in_int[321]), .I (
         uni_cell_in[321])) ;
    IBUF \uni_cell_in_ibuf(322)  (.O (uni_cell_in_int[322]), .I (
         uni_cell_in[322])) ;
    IBUF \uni_cell_in_ibuf(323)  (.O (uni_cell_in_int[323]), .I (
         uni_cell_in[323])) ;
    IBUF \uni_cell_in_ibuf(324)  (.O (uni_cell_in_int[324]), .I (
         uni_cell_in[324])) ;
    IBUF \uni_cell_in_ibuf(325)  (.O (uni_cell_in_int[325]), .I (
         uni_cell_in[325])) ;
    IBUF \uni_cell_in_ibuf(326)  (.O (uni_cell_in_int[326]), .I (
         uni_cell_in[326])) ;
    IBUF \uni_cell_in_ibuf(327)  (.O (uni_cell_in_int[327]), .I (
         uni_cell_in[327])) ;
    IBUF \uni_cell_in_ibuf(328)  (.O (uni_cell_in_int[328]), .I (
         uni_cell_in[328])) ;
    IBUF \uni_cell_in_ibuf(329)  (.O (uni_cell_in_int[329]), .I (
         uni_cell_in[329])) ;
    IBUF \uni_cell_in_ibuf(330)  (.O (uni_cell_in_int[330]), .I (
         uni_cell_in[330])) ;
    IBUF \uni_cell_in_ibuf(331)  (.O (uni_cell_in_int[331]), .I (
         uni_cell_in[331])) ;
    IBUF \uni_cell_in_ibuf(332)  (.O (uni_cell_in_int[332]), .I (
         uni_cell_in[332])) ;
    IBUF \uni_cell_in_ibuf(333)  (.O (uni_cell_in_int[333]), .I (
         uni_cell_in[333])) ;
    IBUF \uni_cell_in_ibuf(334)  (.O (uni_cell_in_int[334]), .I (
         uni_cell_in[334])) ;
    IBUF \uni_cell_in_ibuf(335)  (.O (uni_cell_in_int[335]), .I (
         uni_cell_in[335])) ;
    IBUF \uni_cell_in_ibuf(336)  (.O (uni_cell_in_int[336]), .I (
         uni_cell_in[336])) ;
    IBUF \uni_cell_in_ibuf(337)  (.O (uni_cell_in_int[337]), .I (
         uni_cell_in[337])) ;
    IBUF \uni_cell_in_ibuf(338)  (.O (uni_cell_in_int[338]), .I (
         uni_cell_in[338])) ;
    IBUF \uni_cell_in_ibuf(339)  (.O (uni_cell_in_int[339]), .I (
         uni_cell_in[339])) ;
    IBUF \uni_cell_in_ibuf(340)  (.O (uni_cell_in_int[340]), .I (
         uni_cell_in[340])) ;
    IBUF \uni_cell_in_ibuf(341)  (.O (uni_cell_in_int[341]), .I (
         uni_cell_in[341])) ;
    IBUF \uni_cell_in_ibuf(342)  (.O (uni_cell_in_int[342]), .I (
         uni_cell_in[342])) ;
    IBUF \uni_cell_in_ibuf(343)  (.O (uni_cell_in_int[343]), .I (
         uni_cell_in[343])) ;
    IBUF \uni_cell_in_ibuf(344)  (.O (uni_cell_in_int[344]), .I (
         uni_cell_in[344])) ;
    IBUF \uni_cell_in_ibuf(345)  (.O (uni_cell_in_int[345]), .I (
         uni_cell_in[345])) ;
    IBUF \uni_cell_in_ibuf(346)  (.O (uni_cell_in_int[346]), .I (
         uni_cell_in[346])) ;
    IBUF \uni_cell_in_ibuf(347)  (.O (uni_cell_in_int[347]), .I (
         uni_cell_in[347])) ;
    IBUF \uni_cell_in_ibuf(348)  (.O (uni_cell_in_int[348]), .I (
         uni_cell_in[348])) ;
    IBUF \uni_cell_in_ibuf(349)  (.O (uni_cell_in_int[349]), .I (
         uni_cell_in[349])) ;
    IBUF \uni_cell_in_ibuf(350)  (.O (uni_cell_in_int[350]), .I (
         uni_cell_in[350])) ;
    IBUF \uni_cell_in_ibuf(351)  (.O (uni_cell_in_int[351]), .I (
         uni_cell_in[351])) ;
    IBUF \uni_cell_in_ibuf(352)  (.O (uni_cell_in_int[352]), .I (
         uni_cell_in[352])) ;
    IBUF \uni_cell_in_ibuf(353)  (.O (uni_cell_in_int[353]), .I (
         uni_cell_in[353])) ;
    IBUF \uni_cell_in_ibuf(354)  (.O (uni_cell_in_int[354]), .I (
         uni_cell_in[354])) ;
    IBUF \uni_cell_in_ibuf(355)  (.O (uni_cell_in_int[355]), .I (
         uni_cell_in[355])) ;
    IBUF \uni_cell_in_ibuf(356)  (.O (uni_cell_in_int[356]), .I (
         uni_cell_in[356])) ;
    IBUF \uni_cell_in_ibuf(357)  (.O (uni_cell_in_int[357]), .I (
         uni_cell_in[357])) ;
    IBUF \uni_cell_in_ibuf(358)  (.O (uni_cell_in_int[358]), .I (
         uni_cell_in[358])) ;
    IBUF \uni_cell_in_ibuf(359)  (.O (uni_cell_in_int[359]), .I (
         uni_cell_in[359])) ;
    IBUF \uni_cell_in_ibuf(360)  (.O (uni_cell_in_int[360]), .I (
         uni_cell_in[360])) ;
    IBUF \uni_cell_in_ibuf(361)  (.O (uni_cell_in_int[361]), .I (
         uni_cell_in[361])) ;
    IBUF \uni_cell_in_ibuf(362)  (.O (uni_cell_in_int[362]), .I (
         uni_cell_in[362])) ;
    IBUF \uni_cell_in_ibuf(363)  (.O (uni_cell_in_int[363]), .I (
         uni_cell_in[363])) ;
    IBUF \uni_cell_in_ibuf(364)  (.O (uni_cell_in_int[364]), .I (
         uni_cell_in[364])) ;
    IBUF \uni_cell_in_ibuf(365)  (.O (uni_cell_in_int[365]), .I (
         uni_cell_in[365])) ;
    IBUF \uni_cell_in_ibuf(366)  (.O (uni_cell_in_int[366]), .I (
         uni_cell_in[366])) ;
    IBUF \uni_cell_in_ibuf(367)  (.O (uni_cell_in_int[367]), .I (
         uni_cell_in[367])) ;
    IBUF \uni_cell_in_ibuf(368)  (.O (uni_cell_in_int[368]), .I (
         uni_cell_in[368])) ;
    IBUF \uni_cell_in_ibuf(369)  (.O (uni_cell_in_int[369]), .I (
         uni_cell_in[369])) ;
    IBUF \uni_cell_in_ibuf(370)  (.O (uni_cell_in_int[370]), .I (
         uni_cell_in[370])) ;
    IBUF \uni_cell_in_ibuf(371)  (.O (uni_cell_in_int[371]), .I (
         uni_cell_in[371])) ;
    IBUF \uni_cell_in_ibuf(372)  (.O (uni_cell_in_int[372]), .I (
         uni_cell_in[372])) ;
    IBUF \uni_cell_in_ibuf(373)  (.O (uni_cell_in_int[373]), .I (
         uni_cell_in[373])) ;
    IBUF \uni_cell_in_ibuf(374)  (.O (uni_cell_in_int[374]), .I (
         uni_cell_in[374])) ;
    IBUF \uni_cell_in_ibuf(375)  (.O (uni_cell_in_int[375]), .I (
         uni_cell_in[375])) ;
    IBUF \uni_cell_in_ibuf(376)  (.O (uni_cell_in_int[376]), .I (
         uni_cell_in[376])) ;
    IBUF \uni_cell_in_ibuf(377)  (.O (uni_cell_in_int[377]), .I (
         uni_cell_in[377])) ;
    IBUF \uni_cell_in_ibuf(378)  (.O (uni_cell_in_int[378]), .I (
         uni_cell_in[378])) ;
    IBUF \uni_cell_in_ibuf(379)  (.O (uni_cell_in_int[379]), .I (
         uni_cell_in[379])) ;
    IBUF \uni_cell_in_ibuf(380)  (.O (uni_cell_in_int[380]), .I (
         uni_cell_in[380])) ;
    IBUF \uni_cell_in_ibuf(381)  (.O (uni_cell_in_int[381]), .I (
         uni_cell_in[381])) ;
    IBUF \uni_cell_in_ibuf(382)  (.O (uni_cell_in_int[382]), .I (
         uni_cell_in[382])) ;
    IBUF \uni_cell_in_ibuf(383)  (.O (uni_cell_in_int[383]), .I (
         uni_cell_in[383])) ;
    IBUF \uni_cell_in_ibuf(384)  (.O (uni_cell_in_int[384]), .I (
         uni_cell_in[384])) ;
    IBUF \uni_cell_in_ibuf(385)  (.O (uni_cell_in_int[385]), .I (
         uni_cell_in[385])) ;
    IBUF \uni_cell_in_ibuf(386)  (.O (uni_cell_in_int[386]), .I (
         uni_cell_in[386])) ;
    IBUF \uni_cell_in_ibuf(387)  (.O (uni_cell_in_int[387]), .I (
         uni_cell_in[387])) ;
    IBUF \uni_cell_in_ibuf(388)  (.O (uni_cell_in_int[388]), .I (
         uni_cell_in[388])) ;
    IBUF \uni_cell_in_ibuf(389)  (.O (uni_cell_in_int[389]), .I (
         uni_cell_in[389])) ;
    IBUF \uni_cell_in_ibuf(390)  (.O (uni_cell_in_int[390]), .I (
         uni_cell_in[390])) ;
    IBUF \uni_cell_in_ibuf(391)  (.O (uni_cell_in_int[391]), .I (
         uni_cell_in[391])) ;
    IBUF \uni_cell_in_ibuf(392)  (.O (uni_cell_in_int[392]), .I (
         uni_cell_in[392])) ;
    IBUF \uni_cell_in_ibuf(393)  (.O (uni_cell_in_int[393]), .I (
         uni_cell_in[393])) ;
    IBUF \uni_cell_in_ibuf(394)  (.O (uni_cell_in_int[394]), .I (
         uni_cell_in[394])) ;
    IBUF \uni_cell_in_ibuf(395)  (.O (uni_cell_in_int[395]), .I (
         uni_cell_in[395])) ;
    IBUF \uni_cell_in_ibuf(396)  (.O (uni_cell_in_int[396]), .I (
         uni_cell_in[396])) ;
    IBUF \uni_cell_in_ibuf(397)  (.O (uni_cell_in_int[397]), .I (
         uni_cell_in[397])) ;
    IBUF \uni_cell_in_ibuf(398)  (.O (uni_cell_in_int[398]), .I (
         uni_cell_in[398])) ;
    IBUF \uni_cell_in_ibuf(399)  (.O (uni_cell_in_int[399]), .I (
         uni_cell_in[399])) ;
    IBUF \uni_cell_in_ibuf(400)  (.O (uni_cell_in_int[400]), .I (
         uni_cell_in[400])) ;
    IBUF \uni_cell_in_ibuf(401)  (.O (uni_cell_in_int[401]), .I (
         uni_cell_in[401])) ;
    IBUF \uni_cell_in_ibuf(402)  (.O (uni_cell_in_int[402]), .I (
         uni_cell_in[402])) ;
    IBUF \uni_cell_in_ibuf(403)  (.O (uni_cell_in_int[403]), .I (
         uni_cell_in[403])) ;
    IBUF \uni_cell_in_ibuf(404)  (.O (uni_cell_in_int[404]), .I (
         uni_cell_in[404])) ;
    IBUF \uni_cell_in_ibuf(405)  (.O (uni_cell_in_int[405]), .I (
         uni_cell_in[405])) ;
    IBUF \uni_cell_in_ibuf(406)  (.O (uni_cell_in_int[406]), .I (
         uni_cell_in[406])) ;
    IBUF \uni_cell_in_ibuf(407)  (.O (uni_cell_in_int[407]), .I (
         uni_cell_in[407])) ;
    IBUF \uni_cell_in_ibuf(408)  (.O (uni_cell_in_int[408]), .I (
         uni_cell_in[408])) ;
    IBUF \uni_cell_in_ibuf(409)  (.O (uni_cell_in_int[409]), .I (
         uni_cell_in[409])) ;
    IBUF \uni_cell_in_ibuf(410)  (.O (uni_cell_in_int[410]), .I (
         uni_cell_in[410])) ;
    IBUF \uni_cell_in_ibuf(411)  (.O (uni_cell_in_int[411]), .I (
         uni_cell_in[411])) ;
    IBUF \uni_cell_in_ibuf(412)  (.O (uni_cell_in_int[412]), .I (
         uni_cell_in[412])) ;
    IBUF \uni_cell_in_ibuf(413)  (.O (uni_cell_in_int[413]), .I (
         uni_cell_in[413])) ;
    IBUF \uni_cell_in_ibuf(414)  (.O (uni_cell_in_int[414]), .I (
         uni_cell_in[414])) ;
    IBUF \uni_cell_in_ibuf(415)  (.O (uni_cell_in_int[415]), .I (
         uni_cell_in[415])) ;
    IBUF \uni_cell_in_ibuf(416)  (.O (uni_cell_in_int[416]), .I (
         uni_cell_in[416])) ;
    IBUF \uni_cell_in_ibuf(417)  (.O (uni_cell_in_int[417]), .I (
         uni_cell_in[417])) ;
    IBUF \uni_cell_in_ibuf(418)  (.O (uni_cell_in_int[418]), .I (
         uni_cell_in[418])) ;
    IBUF \uni_cell_in_ibuf(419)  (.O (uni_cell_in_int[419]), .I (
         uni_cell_in[419])) ;
    IBUF \uni_cell_in_ibuf(420)  (.O (uni_cell_in_int[420]), .I (
         uni_cell_in[420])) ;
    IBUF \uni_cell_in_ibuf(421)  (.O (uni_cell_in_int[421]), .I (
         uni_cell_in[421])) ;
    IBUF \uni_cell_in_ibuf(422)  (.O (uni_cell_in_int[422]), .I (
         uni_cell_in[422])) ;
    IBUF \uni_cell_in_ibuf(423)  (.O (uni_cell_in_int[423]), .I (
         uni_cell_in[423])) ;
    IBUF rstN_ibuf (.O (rstN_int), .I (rstN)) ;
    FDC \reg_uni_cell_out_GFC_in(3)  (.Q (uni_cell_out_GFC_in_dup_0[3]), .D (
        uni_cell_in_int[423]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_GFC_in(2)  (.Q (uni_cell_out_GFC_in_dup_0[2]), .D (
        uni_cell_in_int[422]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_GFC_in(1)  (.Q (uni_cell_out_GFC_in_dup_0[1]), .D (
        uni_cell_in_int[421]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_GFC_in(0)  (.Q (uni_cell_out_GFC_in_dup_0[0]), .D (
        uni_cell_in_int[420]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_VPI_in(7)  (.Q (uni_cell_out_VPI_in_dup_0[7]), .D (
        uni_cell_in_int[419]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_VPI_in(6)  (.Q (uni_cell_out_VPI_in_dup_0[6]), .D (
        uni_cell_in_int[418]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_VPI_in(5)  (.Q (uni_cell_out_VPI_in_dup_0[5]), .D (
        uni_cell_in_int[417]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_VPI_in(4)  (.Q (uni_cell_out_VPI_in_dup_0[4]), .D (
        uni_cell_in_int[416]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_VPI_in(3)  (.Q (uni_cell_out_VPI_in_dup_0[3]), .D (
        uni_cell_in_int[415]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_VPI_in(2)  (.Q (uni_cell_out_VPI_in_dup_0[2]), .D (
        uni_cell_in_int[414]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_VPI_in(1)  (.Q (uni_cell_out_VPI_in_dup_0[1]), .D (
        uni_cell_in_int[413]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_VPI_in(0)  (.Q (uni_cell_out_VPI_in_dup_0[0]), .D (
        uni_cell_in_int[412]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_VCI_in(15)  (.Q (uni_cell_out_VCI_in_dup_0[15]), .D (
        uni_cell_in_int[411]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_VCI_in(14)  (.Q (uni_cell_out_VCI_in_dup_0[14]), .D (
        uni_cell_in_int[410]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_VCI_in(13)  (.Q (uni_cell_out_VCI_in_dup_0[13]), .D (
        uni_cell_in_int[409]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_VCI_in(12)  (.Q (uni_cell_out_VCI_in_dup_0[12]), .D (
        uni_cell_in_int[408]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_VCI_in(11)  (.Q (uni_cell_out_VCI_in_dup_0[11]), .D (
        uni_cell_in_int[407]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_VCI_in(10)  (.Q (uni_cell_out_VCI_in_dup_0[10]), .D (
        uni_cell_in_int[406]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_VCI_in(9)  (.Q (uni_cell_out_VCI_in_dup_0[9]), .D (
        uni_cell_in_int[405]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_VCI_in(8)  (.Q (uni_cell_out_VCI_in_dup_0[8]), .D (
        uni_cell_in_int[404]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_VCI_in(7)  (.Q (uni_cell_out_VCI_in_dup_0[7]), .D (
        uni_cell_in_int[403]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_VCI_in(6)  (.Q (uni_cell_out_VCI_in_dup_0[6]), .D (
        uni_cell_in_int[402]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_VCI_in(5)  (.Q (uni_cell_out_VCI_in_dup_0[5]), .D (
        uni_cell_in_int[401]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_VCI_in(4)  (.Q (uni_cell_out_VCI_in_dup_0[4]), .D (
        uni_cell_in_int[400]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_VCI_in(3)  (.Q (uni_cell_out_VCI_in_dup_0[3]), .D (
        uni_cell_in_int[399]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_VCI_in(2)  (.Q (uni_cell_out_VCI_in_dup_0[2]), .D (
        uni_cell_in_int[398]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_VCI_in(1)  (.Q (uni_cell_out_VCI_in_dup_0[1]), .D (
        uni_cell_in_int[397]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_VCI_in(0)  (.Q (uni_cell_out_VCI_in_dup_0[0]), .D (
        uni_cell_in_int[396]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_PTI_in(2)  (.Q (uni_cell_out_PTI_in_dup_0[2]), .D (
        uni_cell_in_int[395]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_PTI_in(1)  (.Q (uni_cell_out_PTI_in_dup_0[1]), .D (
        uni_cell_in_int[394]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_PTI_in(0)  (.Q (uni_cell_out_PTI_in_dup_0[0]), .D (
        uni_cell_in_int[393]), .C (clk_int), .CLR (not_rstN)) ;
    FDC reg_uni_cell_out_CLP_in (.Q (uni_cell_out_CLP_in_dup_0), .D (
        uni_cell_in_int[392]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_HEC_in(7)  (.Q (uni_cell_out_HEC_in_dup_0[7]), .D (
        uni_cell_in_int[391]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_HEC_in(6)  (.Q (uni_cell_out_HEC_in_dup_0[6]), .D (
        uni_cell_in_int[390]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_HEC_in(5)  (.Q (uni_cell_out_HEC_in_dup_0[5]), .D (
        uni_cell_in_int[389]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_HEC_in(4)  (.Q (uni_cell_out_HEC_in_dup_0[4]), .D (
        uni_cell_in_int[388]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_HEC_in(3)  (.Q (uni_cell_out_HEC_in_dup_0[3]), .D (
        uni_cell_in_int[387]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_HEC_in(2)  (.Q (uni_cell_out_HEC_in_dup_0[2]), .D (
        uni_cell_in_int[386]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_HEC_in(1)  (.Q (uni_cell_out_HEC_in_dup_0[1]), .D (
        uni_cell_in_int[385]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_HEC_in(0)  (.Q (uni_cell_out_HEC_in_dup_0[0]), .D (
        uni_cell_in_int[384]), .C (clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(0)(7)  (.Q (
        \uni_cell_out_Payload_in(0)_dup_0(7)  ), .D (uni_cell_in_int[383]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(0)(6)  (.Q (
        \uni_cell_out_Payload_in(0)_dup_0(6)  ), .D (uni_cell_in_int[382]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(0)(5)  (.Q (
        \uni_cell_out_Payload_in(0)_dup_0(5)  ), .D (uni_cell_in_int[381]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(0)(4)  (.Q (
        \uni_cell_out_Payload_in(0)_dup_0(4)  ), .D (uni_cell_in_int[380]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(0)(3)  (.Q (
        \uni_cell_out_Payload_in(0)_dup_0(3)  ), .D (uni_cell_in_int[379]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(0)(2)  (.Q (
        \uni_cell_out_Payload_in(0)_dup_0(2)  ), .D (uni_cell_in_int[378]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(0)(1)  (.Q (
        \uni_cell_out_Payload_in(0)_dup_0(1)  ), .D (uni_cell_in_int[377]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(0)(0)  (.Q (
        \uni_cell_out_Payload_in(0)_dup_0(0)  ), .D (uni_cell_in_int[376]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(1)(7)  (.Q (
        \uni_cell_out_Payload_in(1)_dup_0(7)  ), .D (uni_cell_in_int[375]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(1)(6)  (.Q (
        \uni_cell_out_Payload_in(1)_dup_0(6)  ), .D (uni_cell_in_int[374]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(1)(5)  (.Q (
        \uni_cell_out_Payload_in(1)_dup_0(5)  ), .D (uni_cell_in_int[373]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(1)(4)  (.Q (
        \uni_cell_out_Payload_in(1)_dup_0(4)  ), .D (uni_cell_in_int[372]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(1)(3)  (.Q (
        \uni_cell_out_Payload_in(1)_dup_0(3)  ), .D (uni_cell_in_int[371]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(1)(2)  (.Q (
        \uni_cell_out_Payload_in(1)_dup_0(2)  ), .D (uni_cell_in_int[370]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(1)(1)  (.Q (
        \uni_cell_out_Payload_in(1)_dup_0(1)  ), .D (uni_cell_in_int[369]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(1)(0)  (.Q (
        \uni_cell_out_Payload_in(1)_dup_0(0)  ), .D (uni_cell_in_int[368]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(2)(7)  (.Q (
        \uni_cell_out_Payload_in(2)_dup_0(7)  ), .D (uni_cell_in_int[367]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(2)(6)  (.Q (
        \uni_cell_out_Payload_in(2)_dup_0(6)  ), .D (uni_cell_in_int[366]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(2)(5)  (.Q (
        \uni_cell_out_Payload_in(2)_dup_0(5)  ), .D (uni_cell_in_int[365]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(2)(4)  (.Q (
        \uni_cell_out_Payload_in(2)_dup_0(4)  ), .D (uni_cell_in_int[364]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(2)(3)  (.Q (
        \uni_cell_out_Payload_in(2)_dup_0(3)  ), .D (uni_cell_in_int[363]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(2)(2)  (.Q (
        \uni_cell_out_Payload_in(2)_dup_0(2)  ), .D (uni_cell_in_int[362]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(2)(1)  (.Q (
        \uni_cell_out_Payload_in(2)_dup_0(1)  ), .D (uni_cell_in_int[361]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(2)(0)  (.Q (
        \uni_cell_out_Payload_in(2)_dup_0(0)  ), .D (uni_cell_in_int[360]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(3)(7)  (.Q (
        \uni_cell_out_Payload_in(3)_dup_0(7)  ), .D (uni_cell_in_int[359]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(3)(6)  (.Q (
        \uni_cell_out_Payload_in(3)_dup_0(6)  ), .D (uni_cell_in_int[358]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(3)(5)  (.Q (
        \uni_cell_out_Payload_in(3)_dup_0(5)  ), .D (uni_cell_in_int[357]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(3)(4)  (.Q (
        \uni_cell_out_Payload_in(3)_dup_0(4)  ), .D (uni_cell_in_int[356]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(3)(3)  (.Q (
        \uni_cell_out_Payload_in(3)_dup_0(3)  ), .D (uni_cell_in_int[355]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(3)(2)  (.Q (
        \uni_cell_out_Payload_in(3)_dup_0(2)  ), .D (uni_cell_in_int[354]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(3)(1)  (.Q (
        \uni_cell_out_Payload_in(3)_dup_0(1)  ), .D (uni_cell_in_int[353]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(3)(0)  (.Q (
        \uni_cell_out_Payload_in(3)_dup_0(0)  ), .D (uni_cell_in_int[352]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(4)(7)  (.Q (
        \uni_cell_out_Payload_in(4)_dup_0(7)  ), .D (uni_cell_in_int[351]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(4)(6)  (.Q (
        \uni_cell_out_Payload_in(4)_dup_0(6)  ), .D (uni_cell_in_int[350]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(4)(5)  (.Q (
        \uni_cell_out_Payload_in(4)_dup_0(5)  ), .D (uni_cell_in_int[349]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(4)(4)  (.Q (
        \uni_cell_out_Payload_in(4)_dup_0(4)  ), .D (uni_cell_in_int[348]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(4)(3)  (.Q (
        \uni_cell_out_Payload_in(4)_dup_0(3)  ), .D (uni_cell_in_int[347]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(4)(2)  (.Q (
        \uni_cell_out_Payload_in(4)_dup_0(2)  ), .D (uni_cell_in_int[346]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(4)(1)  (.Q (
        \uni_cell_out_Payload_in(4)_dup_0(1)  ), .D (uni_cell_in_int[345]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(4)(0)  (.Q (
        \uni_cell_out_Payload_in(4)_dup_0(0)  ), .D (uni_cell_in_int[344]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(5)(7)  (.Q (
        \uni_cell_out_Payload_in(5)_dup_0(7)  ), .D (uni_cell_in_int[343]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(5)(6)  (.Q (
        \uni_cell_out_Payload_in(5)_dup_0(6)  ), .D (uni_cell_in_int[342]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(5)(5)  (.Q (
        \uni_cell_out_Payload_in(5)_dup_0(5)  ), .D (uni_cell_in_int[341]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(5)(4)  (.Q (
        \uni_cell_out_Payload_in(5)_dup_0(4)  ), .D (uni_cell_in_int[340]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(5)(3)  (.Q (
        \uni_cell_out_Payload_in(5)_dup_0(3)  ), .D (uni_cell_in_int[339]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(5)(2)  (.Q (
        \uni_cell_out_Payload_in(5)_dup_0(2)  ), .D (uni_cell_in_int[338]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(5)(1)  (.Q (
        \uni_cell_out_Payload_in(5)_dup_0(1)  ), .D (uni_cell_in_int[337]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(5)(0)  (.Q (
        \uni_cell_out_Payload_in(5)_dup_0(0)  ), .D (uni_cell_in_int[336]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(6)(7)  (.Q (
        \uni_cell_out_Payload_in(6)_dup_0(7)  ), .D (uni_cell_in_int[335]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(6)(6)  (.Q (
        \uni_cell_out_Payload_in(6)_dup_0(6)  ), .D (uni_cell_in_int[334]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(6)(5)  (.Q (
        \uni_cell_out_Payload_in(6)_dup_0(5)  ), .D (uni_cell_in_int[333]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(6)(4)  (.Q (
        \uni_cell_out_Payload_in(6)_dup_0(4)  ), .D (uni_cell_in_int[332]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(6)(3)  (.Q (
        \uni_cell_out_Payload_in(6)_dup_0(3)  ), .D (uni_cell_in_int[331]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(6)(2)  (.Q (
        \uni_cell_out_Payload_in(6)_dup_0(2)  ), .D (uni_cell_in_int[330]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(6)(1)  (.Q (
        \uni_cell_out_Payload_in(6)_dup_0(1)  ), .D (uni_cell_in_int[329]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(6)(0)  (.Q (
        \uni_cell_out_Payload_in(6)_dup_0(0)  ), .D (uni_cell_in_int[328]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(7)(7)  (.Q (
        \uni_cell_out_Payload_in(7)_dup_0(7)  ), .D (uni_cell_in_int[327]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(7)(6)  (.Q (
        \uni_cell_out_Payload_in(7)_dup_0(6)  ), .D (uni_cell_in_int[326]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(7)(5)  (.Q (
        \uni_cell_out_Payload_in(7)_dup_0(5)  ), .D (uni_cell_in_int[325]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(7)(4)  (.Q (
        \uni_cell_out_Payload_in(7)_dup_0(4)  ), .D (uni_cell_in_int[324]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(7)(3)  (.Q (
        \uni_cell_out_Payload_in(7)_dup_0(3)  ), .D (uni_cell_in_int[323]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(7)(2)  (.Q (
        \uni_cell_out_Payload_in(7)_dup_0(2)  ), .D (uni_cell_in_int[322]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(7)(1)  (.Q (
        \uni_cell_out_Payload_in(7)_dup_0(1)  ), .D (uni_cell_in_int[321]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(7)(0)  (.Q (
        \uni_cell_out_Payload_in(7)_dup_0(0)  ), .D (uni_cell_in_int[320]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(8)(7)  (.Q (
        \uni_cell_out_Payload_in(8)_dup_0(7)  ), .D (uni_cell_in_int[319]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(8)(6)  (.Q (
        \uni_cell_out_Payload_in(8)_dup_0(6)  ), .D (uni_cell_in_int[318]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(8)(5)  (.Q (
        \uni_cell_out_Payload_in(8)_dup_0(5)  ), .D (uni_cell_in_int[317]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(8)(4)  (.Q (
        \uni_cell_out_Payload_in(8)_dup_0(4)  ), .D (uni_cell_in_int[316]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(8)(3)  (.Q (
        \uni_cell_out_Payload_in(8)_dup_0(3)  ), .D (uni_cell_in_int[315]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(8)(2)  (.Q (
        \uni_cell_out_Payload_in(8)_dup_0(2)  ), .D (uni_cell_in_int[314]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(8)(1)  (.Q (
        \uni_cell_out_Payload_in(8)_dup_0(1)  ), .D (uni_cell_in_int[313]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(8)(0)  (.Q (
        \uni_cell_out_Payload_in(8)_dup_0(0)  ), .D (uni_cell_in_int[312]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(9)(7)  (.Q (
        \uni_cell_out_Payload_in(9)_dup_0(7)  ), .D (uni_cell_in_int[311]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(9)(6)  (.Q (
        \uni_cell_out_Payload_in(9)_dup_0(6)  ), .D (uni_cell_in_int[310]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(9)(5)  (.Q (
        \uni_cell_out_Payload_in(9)_dup_0(5)  ), .D (uni_cell_in_int[309]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(9)(4)  (.Q (
        \uni_cell_out_Payload_in(9)_dup_0(4)  ), .D (uni_cell_in_int[308]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(9)(3)  (.Q (
        \uni_cell_out_Payload_in(9)_dup_0(3)  ), .D (uni_cell_in_int[307]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(9)(2)  (.Q (
        \uni_cell_out_Payload_in(9)_dup_0(2)  ), .D (uni_cell_in_int[306]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(9)(1)  (.Q (
        \uni_cell_out_Payload_in(9)_dup_0(1)  ), .D (uni_cell_in_int[305]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(9)(0)  (.Q (
        \uni_cell_out_Payload_in(9)_dup_0(0)  ), .D (uni_cell_in_int[304]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(10)(7)  (.Q (
        \uni_cell_out_Payload_in(10)_dup_0(7)  ), .D (uni_cell_in_int[303]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(10)(6)  (.Q (
        \uni_cell_out_Payload_in(10)_dup_0(6)  ), .D (uni_cell_in_int[302]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(10)(5)  (.Q (
        \uni_cell_out_Payload_in(10)_dup_0(5)  ), .D (uni_cell_in_int[301]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(10)(4)  (.Q (
        \uni_cell_out_Payload_in(10)_dup_0(4)  ), .D (uni_cell_in_int[300]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(10)(3)  (.Q (
        \uni_cell_out_Payload_in(10)_dup_0(3)  ), .D (uni_cell_in_int[299]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(10)(2)  (.Q (
        \uni_cell_out_Payload_in(10)_dup_0(2)  ), .D (uni_cell_in_int[298]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(10)(1)  (.Q (
        \uni_cell_out_Payload_in(10)_dup_0(1)  ), .D (uni_cell_in_int[297]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(10)(0)  (.Q (
        \uni_cell_out_Payload_in(10)_dup_0(0)  ), .D (uni_cell_in_int[296]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(11)(7)  (.Q (
        \uni_cell_out_Payload_in(11)_dup_0(7)  ), .D (uni_cell_in_int[295]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(11)(6)  (.Q (
        \uni_cell_out_Payload_in(11)_dup_0(6)  ), .D (uni_cell_in_int[294]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(11)(5)  (.Q (
        \uni_cell_out_Payload_in(11)_dup_0(5)  ), .D (uni_cell_in_int[293]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(11)(4)  (.Q (
        \uni_cell_out_Payload_in(11)_dup_0(4)  ), .D (uni_cell_in_int[292]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(11)(3)  (.Q (
        \uni_cell_out_Payload_in(11)_dup_0(3)  ), .D (uni_cell_in_int[291]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(11)(2)  (.Q (
        \uni_cell_out_Payload_in(11)_dup_0(2)  ), .D (uni_cell_in_int[290]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(11)(1)  (.Q (
        \uni_cell_out_Payload_in(11)_dup_0(1)  ), .D (uni_cell_in_int[289]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(11)(0)  (.Q (
        \uni_cell_out_Payload_in(11)_dup_0(0)  ), .D (uni_cell_in_int[288]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(12)(7)  (.Q (
        \uni_cell_out_Payload_in(12)_dup_0(7)  ), .D (uni_cell_in_int[287]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(12)(6)  (.Q (
        \uni_cell_out_Payload_in(12)_dup_0(6)  ), .D (uni_cell_in_int[286]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(12)(5)  (.Q (
        \uni_cell_out_Payload_in(12)_dup_0(5)  ), .D (uni_cell_in_int[285]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(12)(4)  (.Q (
        \uni_cell_out_Payload_in(12)_dup_0(4)  ), .D (uni_cell_in_int[284]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(12)(3)  (.Q (
        \uni_cell_out_Payload_in(12)_dup_0(3)  ), .D (uni_cell_in_int[283]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(12)(2)  (.Q (
        \uni_cell_out_Payload_in(12)_dup_0(2)  ), .D (uni_cell_in_int[282]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(12)(1)  (.Q (
        \uni_cell_out_Payload_in(12)_dup_0(1)  ), .D (uni_cell_in_int[281]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(12)(0)  (.Q (
        \uni_cell_out_Payload_in(12)_dup_0(0)  ), .D (uni_cell_in_int[280]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(13)(7)  (.Q (
        \uni_cell_out_Payload_in(13)_dup_0(7)  ), .D (uni_cell_in_int[279]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(13)(6)  (.Q (
        \uni_cell_out_Payload_in(13)_dup_0(6)  ), .D (uni_cell_in_int[278]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(13)(5)  (.Q (
        \uni_cell_out_Payload_in(13)_dup_0(5)  ), .D (uni_cell_in_int[277]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(13)(4)  (.Q (
        \uni_cell_out_Payload_in(13)_dup_0(4)  ), .D (uni_cell_in_int[276]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(13)(3)  (.Q (
        \uni_cell_out_Payload_in(13)_dup_0(3)  ), .D (uni_cell_in_int[275]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(13)(2)  (.Q (
        \uni_cell_out_Payload_in(13)_dup_0(2)  ), .D (uni_cell_in_int[274]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(13)(1)  (.Q (
        \uni_cell_out_Payload_in(13)_dup_0(1)  ), .D (uni_cell_in_int[273]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(13)(0)  (.Q (
        \uni_cell_out_Payload_in(13)_dup_0(0)  ), .D (uni_cell_in_int[272]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(14)(7)  (.Q (
        \uni_cell_out_Payload_in(14)_dup_0(7)  ), .D (uni_cell_in_int[271]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(14)(6)  (.Q (
        \uni_cell_out_Payload_in(14)_dup_0(6)  ), .D (uni_cell_in_int[270]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(14)(5)  (.Q (
        \uni_cell_out_Payload_in(14)_dup_0(5)  ), .D (uni_cell_in_int[269]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(14)(4)  (.Q (
        \uni_cell_out_Payload_in(14)_dup_0(4)  ), .D (uni_cell_in_int[268]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(14)(3)  (.Q (
        \uni_cell_out_Payload_in(14)_dup_0(3)  ), .D (uni_cell_in_int[267]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(14)(2)  (.Q (
        \uni_cell_out_Payload_in(14)_dup_0(2)  ), .D (uni_cell_in_int[266]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(14)(1)  (.Q (
        \uni_cell_out_Payload_in(14)_dup_0(1)  ), .D (uni_cell_in_int[265]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(14)(0)  (.Q (
        \uni_cell_out_Payload_in(14)_dup_0(0)  ), .D (uni_cell_in_int[264]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(15)(7)  (.Q (
        \uni_cell_out_Payload_in(15)_dup_0(7)  ), .D (uni_cell_in_int[263]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(15)(6)  (.Q (
        \uni_cell_out_Payload_in(15)_dup_0(6)  ), .D (uni_cell_in_int[262]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(15)(5)  (.Q (
        \uni_cell_out_Payload_in(15)_dup_0(5)  ), .D (uni_cell_in_int[261]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(15)(4)  (.Q (
        \uni_cell_out_Payload_in(15)_dup_0(4)  ), .D (uni_cell_in_int[260]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(15)(3)  (.Q (
        \uni_cell_out_Payload_in(15)_dup_0(3)  ), .D (uni_cell_in_int[259]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(15)(2)  (.Q (
        \uni_cell_out_Payload_in(15)_dup_0(2)  ), .D (uni_cell_in_int[258]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(15)(1)  (.Q (
        \uni_cell_out_Payload_in(15)_dup_0(1)  ), .D (uni_cell_in_int[257]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(15)(0)  (.Q (
        \uni_cell_out_Payload_in(15)_dup_0(0)  ), .D (uni_cell_in_int[256]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(16)(7)  (.Q (
        \uni_cell_out_Payload_in(16)_dup_0(7)  ), .D (uni_cell_in_int[255]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(16)(6)  (.Q (
        \uni_cell_out_Payload_in(16)_dup_0(6)  ), .D (uni_cell_in_int[254]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(16)(5)  (.Q (
        \uni_cell_out_Payload_in(16)_dup_0(5)  ), .D (uni_cell_in_int[253]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(16)(4)  (.Q (
        \uni_cell_out_Payload_in(16)_dup_0(4)  ), .D (uni_cell_in_int[252]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(16)(3)  (.Q (
        \uni_cell_out_Payload_in(16)_dup_0(3)  ), .D (uni_cell_in_int[251]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(16)(2)  (.Q (
        \uni_cell_out_Payload_in(16)_dup_0(2)  ), .D (uni_cell_in_int[250]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(16)(1)  (.Q (
        \uni_cell_out_Payload_in(16)_dup_0(1)  ), .D (uni_cell_in_int[249]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(16)(0)  (.Q (
        \uni_cell_out_Payload_in(16)_dup_0(0)  ), .D (uni_cell_in_int[248]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(17)(7)  (.Q (
        \uni_cell_out_Payload_in(17)_dup_0(7)  ), .D (uni_cell_in_int[247]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(17)(6)  (.Q (
        \uni_cell_out_Payload_in(17)_dup_0(6)  ), .D (uni_cell_in_int[246]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(17)(5)  (.Q (
        \uni_cell_out_Payload_in(17)_dup_0(5)  ), .D (uni_cell_in_int[245]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(17)(4)  (.Q (
        \uni_cell_out_Payload_in(17)_dup_0(4)  ), .D (uni_cell_in_int[244]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(17)(3)  (.Q (
        \uni_cell_out_Payload_in(17)_dup_0(3)  ), .D (uni_cell_in_int[243]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(17)(2)  (.Q (
        \uni_cell_out_Payload_in(17)_dup_0(2)  ), .D (uni_cell_in_int[242]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(17)(1)  (.Q (
        \uni_cell_out_Payload_in(17)_dup_0(1)  ), .D (uni_cell_in_int[241]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(17)(0)  (.Q (
        \uni_cell_out_Payload_in(17)_dup_0(0)  ), .D (uni_cell_in_int[240]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(18)(7)  (.Q (
        \uni_cell_out_Payload_in(18)_dup_0(7)  ), .D (uni_cell_in_int[239]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(18)(6)  (.Q (
        \uni_cell_out_Payload_in(18)_dup_0(6)  ), .D (uni_cell_in_int[238]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(18)(5)  (.Q (
        \uni_cell_out_Payload_in(18)_dup_0(5)  ), .D (uni_cell_in_int[237]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(18)(4)  (.Q (
        \uni_cell_out_Payload_in(18)_dup_0(4)  ), .D (uni_cell_in_int[236]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(18)(3)  (.Q (
        \uni_cell_out_Payload_in(18)_dup_0(3)  ), .D (uni_cell_in_int[235]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(18)(2)  (.Q (
        \uni_cell_out_Payload_in(18)_dup_0(2)  ), .D (uni_cell_in_int[234]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(18)(1)  (.Q (
        \uni_cell_out_Payload_in(18)_dup_0(1)  ), .D (uni_cell_in_int[233]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(18)(0)  (.Q (
        \uni_cell_out_Payload_in(18)_dup_0(0)  ), .D (uni_cell_in_int[232]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(19)(7)  (.Q (
        \uni_cell_out_Payload_in(19)_dup_0(7)  ), .D (uni_cell_in_int[231]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(19)(6)  (.Q (
        \uni_cell_out_Payload_in(19)_dup_0(6)  ), .D (uni_cell_in_int[230]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(19)(5)  (.Q (
        \uni_cell_out_Payload_in(19)_dup_0(5)  ), .D (uni_cell_in_int[229]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(19)(4)  (.Q (
        \uni_cell_out_Payload_in(19)_dup_0(4)  ), .D (uni_cell_in_int[228]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(19)(3)  (.Q (
        \uni_cell_out_Payload_in(19)_dup_0(3)  ), .D (uni_cell_in_int[227]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(19)(2)  (.Q (
        \uni_cell_out_Payload_in(19)_dup_0(2)  ), .D (uni_cell_in_int[226]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(19)(1)  (.Q (
        \uni_cell_out_Payload_in(19)_dup_0(1)  ), .D (uni_cell_in_int[225]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(19)(0)  (.Q (
        \uni_cell_out_Payload_in(19)_dup_0(0)  ), .D (uni_cell_in_int[224]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(20)(7)  (.Q (
        \uni_cell_out_Payload_in(20)_dup_0(7)  ), .D (uni_cell_in_int[223]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(20)(6)  (.Q (
        \uni_cell_out_Payload_in(20)_dup_0(6)  ), .D (uni_cell_in_int[222]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(20)(5)  (.Q (
        \uni_cell_out_Payload_in(20)_dup_0(5)  ), .D (uni_cell_in_int[221]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(20)(4)  (.Q (
        \uni_cell_out_Payload_in(20)_dup_0(4)  ), .D (uni_cell_in_int[220]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(20)(3)  (.Q (
        \uni_cell_out_Payload_in(20)_dup_0(3)  ), .D (uni_cell_in_int[219]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(20)(2)  (.Q (
        \uni_cell_out_Payload_in(20)_dup_0(2)  ), .D (uni_cell_in_int[218]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(20)(1)  (.Q (
        \uni_cell_out_Payload_in(20)_dup_0(1)  ), .D (uni_cell_in_int[217]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(20)(0)  (.Q (
        \uni_cell_out_Payload_in(20)_dup_0(0)  ), .D (uni_cell_in_int[216]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(21)(7)  (.Q (
        \uni_cell_out_Payload_in(21)_dup_0(7)  ), .D (uni_cell_in_int[215]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(21)(6)  (.Q (
        \uni_cell_out_Payload_in(21)_dup_0(6)  ), .D (uni_cell_in_int[214]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(21)(5)  (.Q (
        \uni_cell_out_Payload_in(21)_dup_0(5)  ), .D (uni_cell_in_int[213]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(21)(4)  (.Q (
        \uni_cell_out_Payload_in(21)_dup_0(4)  ), .D (uni_cell_in_int[212]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(21)(3)  (.Q (
        \uni_cell_out_Payload_in(21)_dup_0(3)  ), .D (uni_cell_in_int[211]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(21)(2)  (.Q (
        \uni_cell_out_Payload_in(21)_dup_0(2)  ), .D (uni_cell_in_int[210]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(21)(1)  (.Q (
        \uni_cell_out_Payload_in(21)_dup_0(1)  ), .D (uni_cell_in_int[209]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(21)(0)  (.Q (
        \uni_cell_out_Payload_in(21)_dup_0(0)  ), .D (uni_cell_in_int[208]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(22)(7)  (.Q (
        \uni_cell_out_Payload_in(22)_dup_0(7)  ), .D (uni_cell_in_int[207]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(22)(6)  (.Q (
        \uni_cell_out_Payload_in(22)_dup_0(6)  ), .D (uni_cell_in_int[206]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(22)(5)  (.Q (
        \uni_cell_out_Payload_in(22)_dup_0(5)  ), .D (uni_cell_in_int[205]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(22)(4)  (.Q (
        \uni_cell_out_Payload_in(22)_dup_0(4)  ), .D (uni_cell_in_int[204]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(22)(3)  (.Q (
        \uni_cell_out_Payload_in(22)_dup_0(3)  ), .D (uni_cell_in_int[203]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(22)(2)  (.Q (
        \uni_cell_out_Payload_in(22)_dup_0(2)  ), .D (uni_cell_in_int[202]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(22)(1)  (.Q (
        \uni_cell_out_Payload_in(22)_dup_0(1)  ), .D (uni_cell_in_int[201]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(22)(0)  (.Q (
        \uni_cell_out_Payload_in(22)_dup_0(0)  ), .D (uni_cell_in_int[200]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(23)(7)  (.Q (
        \uni_cell_out_Payload_in(23)_dup_0(7)  ), .D (uni_cell_in_int[199]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(23)(6)  (.Q (
        \uni_cell_out_Payload_in(23)_dup_0(6)  ), .D (uni_cell_in_int[198]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(23)(5)  (.Q (
        \uni_cell_out_Payload_in(23)_dup_0(5)  ), .D (uni_cell_in_int[197]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(23)(4)  (.Q (
        \uni_cell_out_Payload_in(23)_dup_0(4)  ), .D (uni_cell_in_int[196]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(23)(3)  (.Q (
        \uni_cell_out_Payload_in(23)_dup_0(3)  ), .D (uni_cell_in_int[195]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(23)(2)  (.Q (
        \uni_cell_out_Payload_in(23)_dup_0(2)  ), .D (uni_cell_in_int[194]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(23)(1)  (.Q (
        \uni_cell_out_Payload_in(23)_dup_0(1)  ), .D (uni_cell_in_int[193]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(23)(0)  (.Q (
        \uni_cell_out_Payload_in(23)_dup_0(0)  ), .D (uni_cell_in_int[192]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(24)(7)  (.Q (
        \uni_cell_out_Payload_in(24)_dup_0(7)  ), .D (uni_cell_in_int[191]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(24)(6)  (.Q (
        \uni_cell_out_Payload_in(24)_dup_0(6)  ), .D (uni_cell_in_int[190]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(24)(5)  (.Q (
        \uni_cell_out_Payload_in(24)_dup_0(5)  ), .D (uni_cell_in_int[189]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(24)(4)  (.Q (
        \uni_cell_out_Payload_in(24)_dup_0(4)  ), .D (uni_cell_in_int[188]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(24)(3)  (.Q (
        \uni_cell_out_Payload_in(24)_dup_0(3)  ), .D (uni_cell_in_int[187]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(24)(2)  (.Q (
        \uni_cell_out_Payload_in(24)_dup_0(2)  ), .D (uni_cell_in_int[186]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(24)(1)  (.Q (
        \uni_cell_out_Payload_in(24)_dup_0(1)  ), .D (uni_cell_in_int[185]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(24)(0)  (.Q (
        \uni_cell_out_Payload_in(24)_dup_0(0)  ), .D (uni_cell_in_int[184]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(25)(7)  (.Q (
        \uni_cell_out_Payload_in(25)_dup_0(7)  ), .D (uni_cell_in_int[183]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(25)(6)  (.Q (
        \uni_cell_out_Payload_in(25)_dup_0(6)  ), .D (uni_cell_in_int[182]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(25)(5)  (.Q (
        \uni_cell_out_Payload_in(25)_dup_0(5)  ), .D (uni_cell_in_int[181]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(25)(4)  (.Q (
        \uni_cell_out_Payload_in(25)_dup_0(4)  ), .D (uni_cell_in_int[180]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(25)(3)  (.Q (
        \uni_cell_out_Payload_in(25)_dup_0(3)  ), .D (uni_cell_in_int[179]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(25)(2)  (.Q (
        \uni_cell_out_Payload_in(25)_dup_0(2)  ), .D (uni_cell_in_int[178]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(25)(1)  (.Q (
        \uni_cell_out_Payload_in(25)_dup_0(1)  ), .D (uni_cell_in_int[177]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(25)(0)  (.Q (
        \uni_cell_out_Payload_in(25)_dup_0(0)  ), .D (uni_cell_in_int[176]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(26)(7)  (.Q (
        \uni_cell_out_Payload_in(26)_dup_0(7)  ), .D (uni_cell_in_int[175]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(26)(6)  (.Q (
        \uni_cell_out_Payload_in(26)_dup_0(6)  ), .D (uni_cell_in_int[174]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(26)(5)  (.Q (
        \uni_cell_out_Payload_in(26)_dup_0(5)  ), .D (uni_cell_in_int[173]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(26)(4)  (.Q (
        \uni_cell_out_Payload_in(26)_dup_0(4)  ), .D (uni_cell_in_int[172]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(26)(3)  (.Q (
        \uni_cell_out_Payload_in(26)_dup_0(3)  ), .D (uni_cell_in_int[171]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(26)(2)  (.Q (
        \uni_cell_out_Payload_in(26)_dup_0(2)  ), .D (uni_cell_in_int[170]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(26)(1)  (.Q (
        \uni_cell_out_Payload_in(26)_dup_0(1)  ), .D (uni_cell_in_int[169]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(26)(0)  (.Q (
        \uni_cell_out_Payload_in(26)_dup_0(0)  ), .D (uni_cell_in_int[168]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(27)(7)  (.Q (
        \uni_cell_out_Payload_in(27)_dup_0(7)  ), .D (uni_cell_in_int[167]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(27)(6)  (.Q (
        \uni_cell_out_Payload_in(27)_dup_0(6)  ), .D (uni_cell_in_int[166]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(27)(5)  (.Q (
        \uni_cell_out_Payload_in(27)_dup_0(5)  ), .D (uni_cell_in_int[165]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(27)(4)  (.Q (
        \uni_cell_out_Payload_in(27)_dup_0(4)  ), .D (uni_cell_in_int[164]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(27)(3)  (.Q (
        \uni_cell_out_Payload_in(27)_dup_0(3)  ), .D (uni_cell_in_int[163]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(27)(2)  (.Q (
        \uni_cell_out_Payload_in(27)_dup_0(2)  ), .D (uni_cell_in_int[162]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(27)(1)  (.Q (
        \uni_cell_out_Payload_in(27)_dup_0(1)  ), .D (uni_cell_in_int[161]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(27)(0)  (.Q (
        \uni_cell_out_Payload_in(27)_dup_0(0)  ), .D (uni_cell_in_int[160]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(28)(7)  (.Q (
        \uni_cell_out_Payload_in(28)_dup_0(7)  ), .D (uni_cell_in_int[159]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(28)(6)  (.Q (
        \uni_cell_out_Payload_in(28)_dup_0(6)  ), .D (uni_cell_in_int[158]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(28)(5)  (.Q (
        \uni_cell_out_Payload_in(28)_dup_0(5)  ), .D (uni_cell_in_int[157]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(28)(4)  (.Q (
        \uni_cell_out_Payload_in(28)_dup_0(4)  ), .D (uni_cell_in_int[156]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(28)(3)  (.Q (
        \uni_cell_out_Payload_in(28)_dup_0(3)  ), .D (uni_cell_in_int[155]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(28)(2)  (.Q (
        \uni_cell_out_Payload_in(28)_dup_0(2)  ), .D (uni_cell_in_int[154]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(28)(1)  (.Q (
        \uni_cell_out_Payload_in(28)_dup_0(1)  ), .D (uni_cell_in_int[153]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(28)(0)  (.Q (
        \uni_cell_out_Payload_in(28)_dup_0(0)  ), .D (uni_cell_in_int[152]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(29)(7)  (.Q (
        \uni_cell_out_Payload_in(29)_dup_0(7)  ), .D (uni_cell_in_int[151]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(29)(6)  (.Q (
        \uni_cell_out_Payload_in(29)_dup_0(6)  ), .D (uni_cell_in_int[150]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(29)(5)  (.Q (
        \uni_cell_out_Payload_in(29)_dup_0(5)  ), .D (uni_cell_in_int[149]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(29)(4)  (.Q (
        \uni_cell_out_Payload_in(29)_dup_0(4)  ), .D (uni_cell_in_int[148]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(29)(3)  (.Q (
        \uni_cell_out_Payload_in(29)_dup_0(3)  ), .D (uni_cell_in_int[147]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(29)(2)  (.Q (
        \uni_cell_out_Payload_in(29)_dup_0(2)  ), .D (uni_cell_in_int[146]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(29)(1)  (.Q (
        \uni_cell_out_Payload_in(29)_dup_0(1)  ), .D (uni_cell_in_int[145]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(29)(0)  (.Q (
        \uni_cell_out_Payload_in(29)_dup_0(0)  ), .D (uni_cell_in_int[144]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(30)(7)  (.Q (
        \uni_cell_out_Payload_in(30)_dup_0(7)  ), .D (uni_cell_in_int[143]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(30)(6)  (.Q (
        \uni_cell_out_Payload_in(30)_dup_0(6)  ), .D (uni_cell_in_int[142]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(30)(5)  (.Q (
        \uni_cell_out_Payload_in(30)_dup_0(5)  ), .D (uni_cell_in_int[141]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(30)(4)  (.Q (
        \uni_cell_out_Payload_in(30)_dup_0(4)  ), .D (uni_cell_in_int[140]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(30)(3)  (.Q (
        \uni_cell_out_Payload_in(30)_dup_0(3)  ), .D (uni_cell_in_int[139]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(30)(2)  (.Q (
        \uni_cell_out_Payload_in(30)_dup_0(2)  ), .D (uni_cell_in_int[138]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(30)(1)  (.Q (
        \uni_cell_out_Payload_in(30)_dup_0(1)  ), .D (uni_cell_in_int[137]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(30)(0)  (.Q (
        \uni_cell_out_Payload_in(30)_dup_0(0)  ), .D (uni_cell_in_int[136]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(31)(7)  (.Q (
        \uni_cell_out_Payload_in(31)_dup_0(7)  ), .D (uni_cell_in_int[135]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(31)(6)  (.Q (
        \uni_cell_out_Payload_in(31)_dup_0(6)  ), .D (uni_cell_in_int[134]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(31)(5)  (.Q (
        \uni_cell_out_Payload_in(31)_dup_0(5)  ), .D (uni_cell_in_int[133]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(31)(4)  (.Q (
        \uni_cell_out_Payload_in(31)_dup_0(4)  ), .D (uni_cell_in_int[132]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(31)(3)  (.Q (
        \uni_cell_out_Payload_in(31)_dup_0(3)  ), .D (uni_cell_in_int[131]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(31)(2)  (.Q (
        \uni_cell_out_Payload_in(31)_dup_0(2)  ), .D (uni_cell_in_int[130]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(31)(1)  (.Q (
        \uni_cell_out_Payload_in(31)_dup_0(1)  ), .D (uni_cell_in_int[129]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(31)(0)  (.Q (
        \uni_cell_out_Payload_in(31)_dup_0(0)  ), .D (uni_cell_in_int[128]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(32)(7)  (.Q (
        \uni_cell_out_Payload_in(32)_dup_0(7)  ), .D (uni_cell_in_int[127]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(32)(6)  (.Q (
        \uni_cell_out_Payload_in(32)_dup_0(6)  ), .D (uni_cell_in_int[126]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(32)(5)  (.Q (
        \uni_cell_out_Payload_in(32)_dup_0(5)  ), .D (uni_cell_in_int[125]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(32)(4)  (.Q (
        \uni_cell_out_Payload_in(32)_dup_0(4)  ), .D (uni_cell_in_int[124]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(32)(3)  (.Q (
        \uni_cell_out_Payload_in(32)_dup_0(3)  ), .D (uni_cell_in_int[123]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(32)(2)  (.Q (
        \uni_cell_out_Payload_in(32)_dup_0(2)  ), .D (uni_cell_in_int[122]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(32)(1)  (.Q (
        \uni_cell_out_Payload_in(32)_dup_0(1)  ), .D (uni_cell_in_int[121]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(32)(0)  (.Q (
        \uni_cell_out_Payload_in(32)_dup_0(0)  ), .D (uni_cell_in_int[120]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(33)(7)  (.Q (
        \uni_cell_out_Payload_in(33)_dup_0(7)  ), .D (uni_cell_in_int[119]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(33)(6)  (.Q (
        \uni_cell_out_Payload_in(33)_dup_0(6)  ), .D (uni_cell_in_int[118]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(33)(5)  (.Q (
        \uni_cell_out_Payload_in(33)_dup_0(5)  ), .D (uni_cell_in_int[117]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(33)(4)  (.Q (
        \uni_cell_out_Payload_in(33)_dup_0(4)  ), .D (uni_cell_in_int[116]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(33)(3)  (.Q (
        \uni_cell_out_Payload_in(33)_dup_0(3)  ), .D (uni_cell_in_int[115]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(33)(2)  (.Q (
        \uni_cell_out_Payload_in(33)_dup_0(2)  ), .D (uni_cell_in_int[114]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(33)(1)  (.Q (
        \uni_cell_out_Payload_in(33)_dup_0(1)  ), .D (uni_cell_in_int[113]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(33)(0)  (.Q (
        \uni_cell_out_Payload_in(33)_dup_0(0)  ), .D (uni_cell_in_int[112]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(34)(7)  (.Q (
        \uni_cell_out_Payload_in(34)_dup_0(7)  ), .D (uni_cell_in_int[111]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(34)(6)  (.Q (
        \uni_cell_out_Payload_in(34)_dup_0(6)  ), .D (uni_cell_in_int[110]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(34)(5)  (.Q (
        \uni_cell_out_Payload_in(34)_dup_0(5)  ), .D (uni_cell_in_int[109]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(34)(4)  (.Q (
        \uni_cell_out_Payload_in(34)_dup_0(4)  ), .D (uni_cell_in_int[108]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(34)(3)  (.Q (
        \uni_cell_out_Payload_in(34)_dup_0(3)  ), .D (uni_cell_in_int[107]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(34)(2)  (.Q (
        \uni_cell_out_Payload_in(34)_dup_0(2)  ), .D (uni_cell_in_int[106]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(34)(1)  (.Q (
        \uni_cell_out_Payload_in(34)_dup_0(1)  ), .D (uni_cell_in_int[105]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(34)(0)  (.Q (
        \uni_cell_out_Payload_in(34)_dup_0(0)  ), .D (uni_cell_in_int[104]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(35)(7)  (.Q (
        \uni_cell_out_Payload_in(35)_dup_0(7)  ), .D (uni_cell_in_int[103]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(35)(6)  (.Q (
        \uni_cell_out_Payload_in(35)_dup_0(6)  ), .D (uni_cell_in_int[102]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(35)(5)  (.Q (
        \uni_cell_out_Payload_in(35)_dup_0(5)  ), .D (uni_cell_in_int[101]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(35)(4)  (.Q (
        \uni_cell_out_Payload_in(35)_dup_0(4)  ), .D (uni_cell_in_int[100]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(35)(3)  (.Q (
        \uni_cell_out_Payload_in(35)_dup_0(3)  ), .D (uni_cell_in_int[99]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(35)(2)  (.Q (
        \uni_cell_out_Payload_in(35)_dup_0(2)  ), .D (uni_cell_in_int[98]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(35)(1)  (.Q (
        \uni_cell_out_Payload_in(35)_dup_0(1)  ), .D (uni_cell_in_int[97]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(35)(0)  (.Q (
        \uni_cell_out_Payload_in(35)_dup_0(0)  ), .D (uni_cell_in_int[96]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(36)(7)  (.Q (
        \uni_cell_out_Payload_in(36)_dup_0(7)  ), .D (uni_cell_in_int[95]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(36)(6)  (.Q (
        \uni_cell_out_Payload_in(36)_dup_0(6)  ), .D (uni_cell_in_int[94]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(36)(5)  (.Q (
        \uni_cell_out_Payload_in(36)_dup_0(5)  ), .D (uni_cell_in_int[93]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(36)(4)  (.Q (
        \uni_cell_out_Payload_in(36)_dup_0(4)  ), .D (uni_cell_in_int[92]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(36)(3)  (.Q (
        \uni_cell_out_Payload_in(36)_dup_0(3)  ), .D (uni_cell_in_int[91]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(36)(2)  (.Q (
        \uni_cell_out_Payload_in(36)_dup_0(2)  ), .D (uni_cell_in_int[90]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(36)(1)  (.Q (
        \uni_cell_out_Payload_in(36)_dup_0(1)  ), .D (uni_cell_in_int[89]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(36)(0)  (.Q (
        \uni_cell_out_Payload_in(36)_dup_0(0)  ), .D (uni_cell_in_int[88]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(37)(7)  (.Q (
        \uni_cell_out_Payload_in(37)_dup_0(7)  ), .D (uni_cell_in_int[87]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(37)(6)  (.Q (
        \uni_cell_out_Payload_in(37)_dup_0(6)  ), .D (uni_cell_in_int[86]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(37)(5)  (.Q (
        \uni_cell_out_Payload_in(37)_dup_0(5)  ), .D (uni_cell_in_int[85]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(37)(4)  (.Q (
        \uni_cell_out_Payload_in(37)_dup_0(4)  ), .D (uni_cell_in_int[84]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(37)(3)  (.Q (
        \uni_cell_out_Payload_in(37)_dup_0(3)  ), .D (uni_cell_in_int[83]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(37)(2)  (.Q (
        \uni_cell_out_Payload_in(37)_dup_0(2)  ), .D (uni_cell_in_int[82]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(37)(1)  (.Q (
        \uni_cell_out_Payload_in(37)_dup_0(1)  ), .D (uni_cell_in_int[81]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(37)(0)  (.Q (
        \uni_cell_out_Payload_in(37)_dup_0(0)  ), .D (uni_cell_in_int[80]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(38)(7)  (.Q (
        \uni_cell_out_Payload_in(38)_dup_0(7)  ), .D (uni_cell_in_int[79]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(38)(6)  (.Q (
        \uni_cell_out_Payload_in(38)_dup_0(6)  ), .D (uni_cell_in_int[78]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(38)(5)  (.Q (
        \uni_cell_out_Payload_in(38)_dup_0(5)  ), .D (uni_cell_in_int[77]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(38)(4)  (.Q (
        \uni_cell_out_Payload_in(38)_dup_0(4)  ), .D (uni_cell_in_int[76]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(38)(3)  (.Q (
        \uni_cell_out_Payload_in(38)_dup_0(3)  ), .D (uni_cell_in_int[75]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(38)(2)  (.Q (
        \uni_cell_out_Payload_in(38)_dup_0(2)  ), .D (uni_cell_in_int[74]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(38)(1)  (.Q (
        \uni_cell_out_Payload_in(38)_dup_0(1)  ), .D (uni_cell_in_int[73]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(38)(0)  (.Q (
        \uni_cell_out_Payload_in(38)_dup_0(0)  ), .D (uni_cell_in_int[72]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(39)(7)  (.Q (
        \uni_cell_out_Payload_in(39)_dup_0(7)  ), .D (uni_cell_in_int[71]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(39)(6)  (.Q (
        \uni_cell_out_Payload_in(39)_dup_0(6)  ), .D (uni_cell_in_int[70]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(39)(5)  (.Q (
        \uni_cell_out_Payload_in(39)_dup_0(5)  ), .D (uni_cell_in_int[69]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(39)(4)  (.Q (
        \uni_cell_out_Payload_in(39)_dup_0(4)  ), .D (uni_cell_in_int[68]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(39)(3)  (.Q (
        \uni_cell_out_Payload_in(39)_dup_0(3)  ), .D (uni_cell_in_int[67]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(39)(2)  (.Q (
        \uni_cell_out_Payload_in(39)_dup_0(2)  ), .D (uni_cell_in_int[66]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(39)(1)  (.Q (
        \uni_cell_out_Payload_in(39)_dup_0(1)  ), .D (uni_cell_in_int[65]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(39)(0)  (.Q (
        \uni_cell_out_Payload_in(39)_dup_0(0)  ), .D (uni_cell_in_int[64]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(40)(7)  (.Q (
        \uni_cell_out_Payload_in(40)_dup_0(7)  ), .D (uni_cell_in_int[63]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(40)(6)  (.Q (
        \uni_cell_out_Payload_in(40)_dup_0(6)  ), .D (uni_cell_in_int[62]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(40)(5)  (.Q (
        \uni_cell_out_Payload_in(40)_dup_0(5)  ), .D (uni_cell_in_int[61]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(40)(4)  (.Q (
        \uni_cell_out_Payload_in(40)_dup_0(4)  ), .D (uni_cell_in_int[60]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(40)(3)  (.Q (
        \uni_cell_out_Payload_in(40)_dup_0(3)  ), .D (uni_cell_in_int[59]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(40)(2)  (.Q (
        \uni_cell_out_Payload_in(40)_dup_0(2)  ), .D (uni_cell_in_int[58]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(40)(1)  (.Q (
        \uni_cell_out_Payload_in(40)_dup_0(1)  ), .D (uni_cell_in_int[57]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(40)(0)  (.Q (
        \uni_cell_out_Payload_in(40)_dup_0(0)  ), .D (uni_cell_in_int[56]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(41)(7)  (.Q (
        \uni_cell_out_Payload_in(41)_dup_0(7)  ), .D (uni_cell_in_int[55]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(41)(6)  (.Q (
        \uni_cell_out_Payload_in(41)_dup_0(6)  ), .D (uni_cell_in_int[54]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(41)(5)  (.Q (
        \uni_cell_out_Payload_in(41)_dup_0(5)  ), .D (uni_cell_in_int[53]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(41)(4)  (.Q (
        \uni_cell_out_Payload_in(41)_dup_0(4)  ), .D (uni_cell_in_int[52]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(41)(3)  (.Q (
        \uni_cell_out_Payload_in(41)_dup_0(3)  ), .D (uni_cell_in_int[51]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(41)(2)  (.Q (
        \uni_cell_out_Payload_in(41)_dup_0(2)  ), .D (uni_cell_in_int[50]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(41)(1)  (.Q (
        \uni_cell_out_Payload_in(41)_dup_0(1)  ), .D (uni_cell_in_int[49]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(41)(0)  (.Q (
        \uni_cell_out_Payload_in(41)_dup_0(0)  ), .D (uni_cell_in_int[48]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(42)(7)  (.Q (
        \uni_cell_out_Payload_in(42)_dup_0(7)  ), .D (uni_cell_in_int[47]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(42)(6)  (.Q (
        \uni_cell_out_Payload_in(42)_dup_0(6)  ), .D (uni_cell_in_int[46]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(42)(5)  (.Q (
        \uni_cell_out_Payload_in(42)_dup_0(5)  ), .D (uni_cell_in_int[45]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(42)(4)  (.Q (
        \uni_cell_out_Payload_in(42)_dup_0(4)  ), .D (uni_cell_in_int[44]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(42)(3)  (.Q (
        \uni_cell_out_Payload_in(42)_dup_0(3)  ), .D (uni_cell_in_int[43]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(42)(2)  (.Q (
        \uni_cell_out_Payload_in(42)_dup_0(2)  ), .D (uni_cell_in_int[42]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(42)(1)  (.Q (
        \uni_cell_out_Payload_in(42)_dup_0(1)  ), .D (uni_cell_in_int[41]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(42)(0)  (.Q (
        \uni_cell_out_Payload_in(42)_dup_0(0)  ), .D (uni_cell_in_int[40]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(43)(7)  (.Q (
        \uni_cell_out_Payload_in(43)_dup_0(7)  ), .D (uni_cell_in_int[39]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(43)(6)  (.Q (
        \uni_cell_out_Payload_in(43)_dup_0(6)  ), .D (uni_cell_in_int[38]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(43)(5)  (.Q (
        \uni_cell_out_Payload_in(43)_dup_0(5)  ), .D (uni_cell_in_int[37]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(43)(4)  (.Q (
        \uni_cell_out_Payload_in(43)_dup_0(4)  ), .D (uni_cell_in_int[36]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(43)(3)  (.Q (
        \uni_cell_out_Payload_in(43)_dup_0(3)  ), .D (uni_cell_in_int[35]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(43)(2)  (.Q (
        \uni_cell_out_Payload_in(43)_dup_0(2)  ), .D (uni_cell_in_int[34]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(43)(1)  (.Q (
        \uni_cell_out_Payload_in(43)_dup_0(1)  ), .D (uni_cell_in_int[33]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(43)(0)  (.Q (
        \uni_cell_out_Payload_in(43)_dup_0(0)  ), .D (uni_cell_in_int[32]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(44)(7)  (.Q (
        \uni_cell_out_Payload_in(44)_dup_0(7)  ), .D (uni_cell_in_int[31]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(44)(6)  (.Q (
        \uni_cell_out_Payload_in(44)_dup_0(6)  ), .D (uni_cell_in_int[30]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(44)(5)  (.Q (
        \uni_cell_out_Payload_in(44)_dup_0(5)  ), .D (uni_cell_in_int[29]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(44)(4)  (.Q (
        \uni_cell_out_Payload_in(44)_dup_0(4)  ), .D (uni_cell_in_int[28]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(44)(3)  (.Q (
        \uni_cell_out_Payload_in(44)_dup_0(3)  ), .D (uni_cell_in_int[27]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(44)(2)  (.Q (
        \uni_cell_out_Payload_in(44)_dup_0(2)  ), .D (uni_cell_in_int[26]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(44)(1)  (.Q (
        \uni_cell_out_Payload_in(44)_dup_0(1)  ), .D (uni_cell_in_int[25]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(44)(0)  (.Q (
        \uni_cell_out_Payload_in(44)_dup_0(0)  ), .D (uni_cell_in_int[24]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(45)(7)  (.Q (
        \uni_cell_out_Payload_in(45)_dup_0(7)  ), .D (uni_cell_in_int[23]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(45)(6)  (.Q (
        \uni_cell_out_Payload_in(45)_dup_0(6)  ), .D (uni_cell_in_int[22]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(45)(5)  (.Q (
        \uni_cell_out_Payload_in(45)_dup_0(5)  ), .D (uni_cell_in_int[21]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(45)(4)  (.Q (
        \uni_cell_out_Payload_in(45)_dup_0(4)  ), .D (uni_cell_in_int[20]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(45)(3)  (.Q (
        \uni_cell_out_Payload_in(45)_dup_0(3)  ), .D (uni_cell_in_int[19]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(45)(2)  (.Q (
        \uni_cell_out_Payload_in(45)_dup_0(2)  ), .D (uni_cell_in_int[18]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(45)(1)  (.Q (
        \uni_cell_out_Payload_in(45)_dup_0(1)  ), .D (uni_cell_in_int[17]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(45)(0)  (.Q (
        \uni_cell_out_Payload_in(45)_dup_0(0)  ), .D (uni_cell_in_int[16]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(46)(7)  (.Q (
        \uni_cell_out_Payload_in(46)_dup_0(7)  ), .D (uni_cell_in_int[15]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(46)(6)  (.Q (
        \uni_cell_out_Payload_in(46)_dup_0(6)  ), .D (uni_cell_in_int[14]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(46)(5)  (.Q (
        \uni_cell_out_Payload_in(46)_dup_0(5)  ), .D (uni_cell_in_int[13]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(46)(4)  (.Q (
        \uni_cell_out_Payload_in(46)_dup_0(4)  ), .D (uni_cell_in_int[12]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(46)(3)  (.Q (
        \uni_cell_out_Payload_in(46)_dup_0(3)  ), .D (uni_cell_in_int[11]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(46)(2)  (.Q (
        \uni_cell_out_Payload_in(46)_dup_0(2)  ), .D (uni_cell_in_int[10]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(46)(1)  (.Q (
        \uni_cell_out_Payload_in(46)_dup_0(1)  ), .D (uni_cell_in_int[9]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(46)(0)  (.Q (
        \uni_cell_out_Payload_in(46)_dup_0(0)  ), .D (uni_cell_in_int[8]), .C (
        clk_int), .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(47)(7)  (.Q (
        uni_cell_out_Payload_in_dup_0[7]), .D (uni_cell_in_int[7]), .C (clk_int)
        , .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(47)(6)  (.Q (
        uni_cell_out_Payload_in_dup_0[6]), .D (uni_cell_in_int[6]), .C (clk_int)
        , .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(47)(5)  (.Q (
        uni_cell_out_Payload_in_dup_0[5]), .D (uni_cell_in_int[5]), .C (clk_int)
        , .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(47)(4)  (.Q (
        uni_cell_out_Payload_in_dup_0[4]), .D (uni_cell_in_int[4]), .C (clk_int)
        , .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(47)(3)  (.Q (
        uni_cell_out_Payload_in_dup_0[3]), .D (uni_cell_in_int[3]), .C (clk_int)
        , .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(47)(2)  (.Q (
        uni_cell_out_Payload_in_dup_0[2]), .D (uni_cell_in_int[2]), .C (clk_int)
        , .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(47)(1)  (.Q (
        uni_cell_out_Payload_in_dup_0[1]), .D (uni_cell_in_int[1]), .C (clk_int)
        , .CLR (not_rstN)) ;
    FDC \reg_uni_cell_out_Payload_in(47)(0)  (.Q (
        uni_cell_out_Payload_in_dup_0[0]), .D (uni_cell_in_int[0]), .C (clk_int)
        , .CLR (not_rstN)) ;
    LUT1 ix51434z1315 (.O (not_rstN), .I0 (rstN_int)) ;
         defparam ix51434z1315.INIT = 4'h1;
    BUFGP clk_ibuf (.O (clk_int), .I (clk)) ;
endmodule

