/**********************************************************************
 * Illegal use of variables; SystemVerilog checks that at most one
 * continuous assignment or one output port is "driving" a variable and
 * that a cont. assign or output port is not combined with a procedural
 * assignment to the variable.
 *
 * Author: Stuart Sutherland
 *
 * (c) Copyright 2003, Sutherland HDL, Inc. *** ALL RIGHTS RESERVED ***
 * www.sutherland-hdl.com
 *
 * Used with permission in the book, "SystemVerilog for Design"
 *  By Stuart Sutherland, Simon Davidmann, and Peter Flake.
 *  Book copyright: 2003, Kluwer Academic Publishers, Norwell, MA, USA
 *  www.wkap.il, ISBN: 0-4020-7530-8
 *
 * Revision History:
 *   1.00 15 Dec 2003 -- original code, as included in book
 *   1.01 10 Jul 2004 -- cleaned up comments, added expected results
 *                       to output messages
 *
 * Caveat: Expected results displayed for this code example are based
 * on an interpretation of the SystemVerilog 3.1 standard by the code
 * author or authors.  At the time of writing, official SystemVerilog
 * validation suites were not available to validate the example.
 *
 * RIGHT TO USE: This code example, or any portion thereof, may be
 * used and distributed without restriction, provided that this entire
 * comment block is included with the example.
 *
 * DISCLAIMER: THIS CODE EXAMPLE IS PROVIDED "AS IS" WITHOUT WARRANTY
 * OF ANY KIND, EITHER EXPRESS OR IMPLIED, INCLUDING, BUT NOT LIMITED
 * TO WARRANTIES OF MERCHANTABILITY, FITNESS OR CORRECTNESS. IN NO
 * EVENT SHALL THE AUTHOR OR AUTHORS BE LIABLE FOR ANY DAMAGES,
 * INCLUDING INCIDENTAL OR CONSEQUENTIAL DAMAGES, ARISING OUT OF THE
 * USE OF THIS CODE.
 *********************************************************************/

module add_and_increment (output bit [63:0] sum,
                          output bit        carry,
                          input  bit [63:0] a, b );

  always @(a, b)
    sum = a + b;         // OK: procedural assignment to sum

  assign sum = a + 1;    // ERROR! sum is already being
                            // assigned a value

  look_ahead i1 (carry, a, b);  // module instance drives carry

  overflow_check i2 (carry, a, b); // ERROR! 2nd driver of carry

endmodule

module look_ahead (output wire carry,
                   input  bit [63:0] a, b);
  //...
  assign carry = 1'b0;
endmodule

module overflow_check (output wire carry,
                       input  bit [63:0] a, b);
  //...
  assign carry = 1'b1;
endmodule

module test;
  wire [63:0] sum;
  wire carry;
  bit  [63:0] a, b;

  add_and_increment dut (sum, carry, a, b);

  initial begin
    $display("\nExpect errors regarding multiple sources putting values on sum and carry \n");
    a = 2;
    b = 5;
    #1 $display("\nsum=%0d  carry=%0d (expect compile errors)\n", sum, carry);
    $finish;
  end
endmodule