package router_test_pkg;

import uvm_pkg::*;
import router_stimulus_pkg::*;
import router_env_pkg::*;

`include "test_collection.sv"

endpackage
