//--------------------------------------------------------------------------
// Designer: Macro
// Brief: Direct Cache Design
// Change Log:
//--------------------------------------------------------------------------

//--------------------------------------------------------------------------
// Include File
//--------------------------------------------------------------------------

//--------------------------------------------------------------------------
// Module
//--------------------------------------------------------------------------
module direct_cache
//--------------------------------------------------------------------------
// Params
//--------------------------------------------------------------------------
#(
)
//--------------------------------------------------------------------------
// Ports
//--------------------------------------------------------------------------
(
    // Inputs
    input wire         clk,
    input wire         rst_n, 
    input wire [31:0]  mem_addr


    // Outputs
);


endmodule

//--------------------------------------------------------------------------
