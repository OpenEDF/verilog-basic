//Lab 1 - Task 3, Step 2
//
//Declare a program block with arguments to connect
//to modport TB declared in interface
//ToDo

  //Lab 1 - Task 3, Step 3
  //
  //Declare an initial block 
  //In the initial block print a simple message to the screen
  //ToDo

  //Lab 1 - Task 6, Step 3 
  //
  //Replace $display with a call to the reset() task
  //ToDo - Caution!! Do only in Task 6

  //Lab 1 - Task 6, Step 2
  //
  //Define a task called reset() inside the program to reset DUT per spec.
  //ToDo - Caution!! Do only in Task 6

