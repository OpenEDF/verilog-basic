/**********************************************************************
 * Unpacked array in-line initialization
 *
 * Author: Stuart Sutherland
 *
 * (c) Copyright 2003, Sutherland HDL, Inc. *** ALL RIGHTS RESERVED ***
 * www.sutherland-hdl.com
 *
 * Used with permission in the book, "SystemVerilog for Design"
 *  By Stuart Sutherland, Simon Davidmann, and Peter Flake.
 *  Book copyright: 2003, Kluwer Academic Publishers, Norwell, MA, USA
 *  www.wkap.il, ISBN: 0-4020-7530-8
 *
 * Revision History:
 *   1.00 15 Dec 2003 -- original code, as included in book
 *   1.01 10 Jul 2004 -- cleaned up comments, added expected results
 *                       to output messages
 *
 * Caveat: Expected results displayed for this code example are based
 * on an interpretation of the SystemVerilog 3.1 standard by the code
 * author or authors.  At the time of writing, official SystemVerilog
 * validation suites were not available to validate the example.
 *
 * RIGHT TO USE: This code example, or any portion thereof, may be
 * used and distributed without restriction, provided that this entire
 * comment block is included with the example.
 *
 * DISCLAIMER: THIS CODE EXAMPLE IS PROVIDED "AS IS" WITHOUT WARRANTY
 * OF ANY KIND, EITHER EXPRESS OR IMPLIED, INCLUDING, BUT NOT LIMITED
 * TO WARRANTIES OF MERCHANTABILITY, FITNESS OR CORRECTNESS. IN NO
 * EVENT SHALL THE AUTHOR OR AUTHORS BE LIABLE FOR ANY DAMAGES,
 * INCLUDING INCIDENTAL OR CONSEQUENTIAL DAMAGES, ARISING OUT OF THE
 * USE OF THIS CODE.
 *********************************************************************/

module test;

  int d1 [0:1][0:3] = { {7,3,0,5}, {2,0,1,6} };
  int d2 [0:1][0:3] = { 2{7,3,0,5} };

  initial begin
    $display("\n d1[0][0] = %0d (expect 7)", d1[0][0]);
    $display(" d1[0][1] = %0d (expect 3)", d1[0][1]);
    $display(" d1[0][2] = %0d (expect 0)", d1[0][2]);
    $display(" d1[0][3] = %0d (expect 5)", d1[0][3]);

    $display("\n d1[1][0] = %0d (expect 2)", d1[1][0]);
    $display(" d1[1][1] = %0d (expect 0)", d1[1][1]);
    $display(" d1[1][2] = %0d (expect 1)", d1[1][2]);
    $display(" d1[1][3] = %0d (expect 6)\n)", d1[1][3]);

    $display("\n d2[0][0] = %0d (expect 7)", d2[0][0]);
    $display(" d2[0][1] = %0d (expect 3)", d2[0][1]);
    $display(" d2[0][2] = %0d (expect 0)", d2[0][2]);
    $display(" d2[0][3] = %0d (expect 5)", d2[0][3]);

    $display("\n d2[1][0] = %0d (expect 7)", d2[1][0]);
    $display(" d2[1][1] = %0d (expect 3)", d2[1][1]);
    $display(" d2[1][2] = %0d (expect 0)", d2[1][2]);
    $display(" d2[1][3] = %0d (expect 5)\n)", d2[1][3]);
    $finish;
  end
endmodule
