/* timescale */
`timescale 1ns/10ps

module top (
    input xx,
    input xx,

)
