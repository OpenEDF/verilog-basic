//--------------------------------------------------------------------------
// Designer: Macro
// Brief: Direct Cache Design
// Change Log:
//--------------------------------------------------------------------------

//--------------------------------------------------------------------------
// Include File
//--------------------------------------------------------------------------

//--------------------------------------------------------------------------
// Module
//--------------------------------------------------------------------------
module direct_cache
//--------------------------------------------------------------------------
// Params
//--------------------------------------------------------------------------
#(
    parameter ENTRY = 8,

)
//--------------------------------------------------------------------------
// Ports
//--------------------------------------------------------------------------
(
    // Inputs
    input wire         clk,
    input wire         rst_n, 
    input wire  [31:0] mem_addr

    // Outputs
    output wire        hit,
    output wire [31:0] data
);

// 8 Entry (1+27+32) bit SRAM
reg []

endmodule

//--------------------------------------------------------------------------
